// soc_system_v5.v

// Generated using ACDS version 17.1 590

`timescale 1 ps / 1 ps
module soc_system_v5 (
		input  wire [15:0] adc_fifo_in_data,                          //                 adc_fifo_in.data
		input  wire        adc_fifo_in_valid,                         //                            .valid
		output wire        adc_fifo_in_ready,                         //                            .ready
		output wire [31:0] adc_val_sub_export,                        //                 adc_val_sub.export
		input  wire        alt_vip_itc_0_clocked_video_vid_clk,       // alt_vip_itc_0_clocked_video.vid_clk
		output wire [31:0] alt_vip_itc_0_clocked_video_vid_data,      //                            .vid_data
		output wire        alt_vip_itc_0_clocked_video_underflow,     //                            .underflow
		output wire        alt_vip_itc_0_clocked_video_vid_datavalid, //                            .vid_datavalid
		output wire        alt_vip_itc_0_clocked_video_vid_v_sync,    //                            .vid_v_sync
		output wire        alt_vip_itc_0_clocked_video_vid_h_sync,    //                            .vid_h_sync
		output wire        alt_vip_itc_0_clocked_video_vid_f,         //                            .vid_f
		output wire        alt_vip_itc_0_clocked_video_vid_h,         //                            .vid_h
		output wire        alt_vip_itc_0_clocked_video_vid_v,         //                            .vid_v
		output wire        analyzer_pll_locked_export,                //         analyzer_pll_locked.export
		output wire        analyzer_pll_outclk0_clk,                  //        analyzer_pll_outclk0.clk
		output wire        analyzer_pll_outclk1_clk,                  //        analyzer_pll_outclk1.clk
		output wire        analyzer_pll_outclk2_clk,                  //        analyzer_pll_outclk2.clk
		output wire        analyzer_pll_outclk3_clk,                  //        analyzer_pll_outclk3.clk
		input  wire        analyzer_pll_reset_reset,                  //          analyzer_pll_reset.reset
		output wire [31:0] aux_cnt_out_export,                        //                 aux_cnt_out.export
		input  wire        clk_clk,                                   //                         clk.clk
		input  wire [7:0]  ctrl_in_export,                            //                     ctrl_in.export
		output wire [31:0] ctrl_out_export,                           //                    ctrl_out.export
		input  wire        dac_grad_MISO,                             //                    dac_grad.MISO
		output wire        dac_grad_MOSI,                             //                            .MOSI
		output wire        dac_grad_SCLK,                             //                            .SCLK
		output wire        dac_grad_SS_n,                             //                            .SS_n
		input  wire [31:0] dconv_fifo_in_data,                        //               dconv_fifo_in.data
		input  wire        dconv_fifo_in_valid,                       //                            .valid
		output wire        dconv_fifo_in_ready,                       //                            .ready
		input  wire [31:0] dconv_fifo_q_in_data,                      //             dconv_fifo_q_in.data
		input  wire        dconv_fifo_q_in_valid,                     //                            .valid
		output wire        dconv_fifo_q_in_ready,                     //                            .ready
		input  wire [14:0] dconv_fir_in_data,                         //                dconv_fir_in.data
		input  wire        dconv_fir_in_valid,                        //                            .valid
		input  wire [1:0]  dconv_fir_in_error,                        //                            .error
		output wire [31:0] dconv_fir_out_data,                        //               dconv_fir_out.data
		output wire        dconv_fir_out_valid,                       //                            .valid
		output wire [1:0]  dconv_fir_out_error,                       //                            .error
		input  wire [14:0] dconv_fir_q_in_data,                       //              dconv_fir_q_in.data
		input  wire        dconv_fir_q_in_valid,                      //                            .valid
		input  wire [1:0]  dconv_fir_q_in_error,                      //                            .error
		output wire [31:0] dconv_fir_q_out_data,                      //             dconv_fir_q_out.data
		output wire        dconv_fir_q_out_valid,                     //                            .valid
		output wire [1:0]  dconv_fir_q_out_error,                     //                            .error
		output wire [31:0] delay_nosig_export,                        //                 delay_nosig.export
		output wire [31:0] delay_sig_export,                          //                   delay_sig.export
		output wire [31:0] delay_t1_export,                           //                    delay_t1.export
		output wire [31:0] echoes_per_scan_export,                    //             echoes_per_scan.export
		input  wire        fifo_clk_bridge_in_clk,                    //          fifo_clk_bridge_in.clk
		input  wire        fifo_rst_reset,                            //                    fifo_rst.reset
		output wire        hps_0_h2f_reset_reset_n,                   //             hps_0_h2f_reset.reset_n
		output wire        hps_0_hps_io_hps_io_emac1_inst_TX_CLK,     //                hps_0_hps_io.hps_io_emac1_inst_TX_CLK
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD0,       //                            .hps_io_emac1_inst_TXD0
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD1,       //                            .hps_io_emac1_inst_TXD1
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD2,       //                            .hps_io_emac1_inst_TXD2
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD3,       //                            .hps_io_emac1_inst_TXD3
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD0,       //                            .hps_io_emac1_inst_RXD0
		inout  wire        hps_0_hps_io_hps_io_emac1_inst_MDIO,       //                            .hps_io_emac1_inst_MDIO
		output wire        hps_0_hps_io_hps_io_emac1_inst_MDC,        //                            .hps_io_emac1_inst_MDC
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RX_CTL,     //                            .hps_io_emac1_inst_RX_CTL
		output wire        hps_0_hps_io_hps_io_emac1_inst_TX_CTL,     //                            .hps_io_emac1_inst_TX_CTL
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RX_CLK,     //                            .hps_io_emac1_inst_RX_CLK
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD1,       //                            .hps_io_emac1_inst_RXD1
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD2,       //                            .hps_io_emac1_inst_RXD2
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD3,       //                            .hps_io_emac1_inst_RXD3
		inout  wire        hps_0_hps_io_hps_io_qspi_inst_IO0,         //                            .hps_io_qspi_inst_IO0
		inout  wire        hps_0_hps_io_hps_io_qspi_inst_IO1,         //                            .hps_io_qspi_inst_IO1
		inout  wire        hps_0_hps_io_hps_io_qspi_inst_IO2,         //                            .hps_io_qspi_inst_IO2
		inout  wire        hps_0_hps_io_hps_io_qspi_inst_IO3,         //                            .hps_io_qspi_inst_IO3
		output wire        hps_0_hps_io_hps_io_qspi_inst_SS0,         //                            .hps_io_qspi_inst_SS0
		output wire        hps_0_hps_io_hps_io_qspi_inst_CLK,         //                            .hps_io_qspi_inst_CLK
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_CMD,         //                            .hps_io_sdio_inst_CMD
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D0,          //                            .hps_io_sdio_inst_D0
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D1,          //                            .hps_io_sdio_inst_D1
		output wire        hps_0_hps_io_hps_io_sdio_inst_CLK,         //                            .hps_io_sdio_inst_CLK
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D2,          //                            .hps_io_sdio_inst_D2
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D3,          //                            .hps_io_sdio_inst_D3
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D0,          //                            .hps_io_usb1_inst_D0
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D1,          //                            .hps_io_usb1_inst_D1
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D2,          //                            .hps_io_usb1_inst_D2
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D3,          //                            .hps_io_usb1_inst_D3
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D4,          //                            .hps_io_usb1_inst_D4
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D5,          //                            .hps_io_usb1_inst_D5
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D6,          //                            .hps_io_usb1_inst_D6
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D7,          //                            .hps_io_usb1_inst_D7
		input  wire        hps_0_hps_io_hps_io_usb1_inst_CLK,         //                            .hps_io_usb1_inst_CLK
		output wire        hps_0_hps_io_hps_io_usb1_inst_STP,         //                            .hps_io_usb1_inst_STP
		input  wire        hps_0_hps_io_hps_io_usb1_inst_DIR,         //                            .hps_io_usb1_inst_DIR
		input  wire        hps_0_hps_io_hps_io_usb1_inst_NXT,         //                            .hps_io_usb1_inst_NXT
		output wire        hps_0_hps_io_hps_io_spim1_inst_CLK,        //                            .hps_io_spim1_inst_CLK
		output wire        hps_0_hps_io_hps_io_spim1_inst_MOSI,       //                            .hps_io_spim1_inst_MOSI
		input  wire        hps_0_hps_io_hps_io_spim1_inst_MISO,       //                            .hps_io_spim1_inst_MISO
		output wire        hps_0_hps_io_hps_io_spim1_inst_SS0,        //                            .hps_io_spim1_inst_SS0
		input  wire        hps_0_hps_io_hps_io_uart0_inst_RX,         //                            .hps_io_uart0_inst_RX
		output wire        hps_0_hps_io_hps_io_uart0_inst_TX,         //                            .hps_io_uart0_inst_TX
		inout  wire        hps_0_hps_io_hps_io_i2c0_inst_SDA,         //                            .hps_io_i2c0_inst_SDA
		inout  wire        hps_0_hps_io_hps_io_i2c0_inst_SCL,         //                            .hps_io_i2c0_inst_SCL
		inout  wire        hps_0_hps_io_hps_io_i2c1_inst_SDA,         //                            .hps_io_i2c1_inst_SDA
		inout  wire        hps_0_hps_io_hps_io_i2c1_inst_SCL,         //                            .hps_io_i2c1_inst_SCL
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO09,      //                            .hps_io_gpio_inst_GPIO09
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO35,      //                            .hps_io_gpio_inst_GPIO35
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO40,      //                            .hps_io_gpio_inst_GPIO40
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO48,      //                            .hps_io_gpio_inst_GPIO48
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO53,      //                            .hps_io_gpio_inst_GPIO53
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO54,      //                            .hps_io_gpio_inst_GPIO54
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO61,      //                            .hps_io_gpio_inst_GPIO61
		input  wire        i2c_ext_sda_in,                            //                     i2c_ext.sda_in
		input  wire        i2c_ext_scl_in,                            //                            .scl_in
		output wire        i2c_ext_sda_oe,                            //                            .sda_oe
		output wire        i2c_ext_scl_oe,                            //                            .scl_oe
		input  wire        i2c_int_sda_in,                            //                     i2c_int.sda_in
		input  wire        i2c_int_scl_in,                            //                            .scl_in
		output wire        i2c_int_sda_oe,                            //                            .sda_oe
		output wire        i2c_int_scl_oe,                            //                            .scl_oe
		output wire [31:0] init_delay_export,                         //                  init_delay.export
		output wire [14:0] memory_mem_a,                              //                      memory.mem_a
		output wire [2:0]  memory_mem_ba,                             //                            .mem_ba
		output wire        memory_mem_ck,                             //                            .mem_ck
		output wire        memory_mem_ck_n,                           //                            .mem_ck_n
		output wire        memory_mem_cke,                            //                            .mem_cke
		output wire        memory_mem_cs_n,                           //                            .mem_cs_n
		output wire        memory_mem_ras_n,                          //                            .mem_ras_n
		output wire        memory_mem_cas_n,                          //                            .mem_cas_n
		output wire        memory_mem_we_n,                           //                            .mem_we_n
		output wire        memory_mem_reset_n,                        //                            .mem_reset_n
		inout  wire [31:0] memory_mem_dq,                             //                            .mem_dq
		inout  wire [3:0]  memory_mem_dqs,                            //                            .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,                          //                            .mem_dqs_n
		output wire        memory_mem_odt,                            //                            .mem_odt
		output wire [3:0]  memory_mem_dm,                             //                            .mem_dm
		input  wire        memory_oct_rzqin,                          //                            .oct_rzqin
		output wire        nmr_sys_pll_locked_export,                 //          nmr_sys_pll_locked.export
		output wire        nmr_sys_pll_outclk_clk,                    //          nmr_sys_pll_outclk.clk
		input  wire        nmr_sys_pll_reset_reset,                   //           nmr_sys_pll_reset.reset
		output wire        pll_vga_clk65_clk,                         //               pll_vga_clk65.clk
		output wire        pll_vga_locked_export,                     //              pll_vga_locked.export
		output wire [31:0] pulse_180deg_export,                       //                pulse_180deg.export
		output wire [31:0] pulse_90deg_export,                        //                 pulse_90deg.export
		output wire [31:0] pulse_t1_export,                           //                    pulse_t1.export
		input  wire        reset_reset_n,                             //                       reset.reset_n
		output wire [31:0] rx_delay_export,                           //                    rx_delay.export
		output wire [31:0] samples_per_echo_export,                   //            samples_per_echo.export
		output wire        sdram_clk_clk,                             //                   sdram_clk.clk
		output wire [12:0] sdram_wire_addr,                           //                  sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,                             //                            .ba
		output wire        sdram_wire_cas_n,                          //                            .cas_n
		output wire        sdram_wire_cke,                            //                            .cke
		output wire        sdram_wire_cs_n,                           //                            .cs_n
		inout  wire [15:0] sdram_wire_dq,                             //                            .dq
		output wire [1:0]  sdram_wire_dqm,                            //                            .dqm
		output wire        sdram_wire_ras_n,                          //                            .ras_n
		output wire        sdram_wire_we_n,                           //                            .we_n
		input  wire        spi_afe_relays_MISO,                       //              spi_afe_relays.MISO
		output wire        spi_afe_relays_MOSI,                       //                            .MOSI
		output wire        spi_afe_relays_SCLK,                       //                            .SCLK
		output wire        spi_afe_relays_SS_n,                       //                            .SS_n
		input  wire        spi_mtch_ntwrk_MISO,                       //              spi_mtch_ntwrk.MISO
		output wire        spi_mtch_ntwrk_MOSI,                       //                            .MOSI
		output wire        spi_mtch_ntwrk_SCLK,                       //                            .SCLK
		output wire        spi_mtch_ntwrk_SS_n,                       //                            .SS_n
		input  wire [9:0]  switches_export                            //                    switches.export
	);

	wire          alt_vip_vfr_vga_avalon_streaming_source_valid;                         // alt_vip_vfr_vga:dout_valid -> alt_vip_itc_0:is_valid
	wire   [31:0] alt_vip_vfr_vga_avalon_streaming_source_data;                          // alt_vip_vfr_vga:dout_data -> alt_vip_itc_0:is_data
	wire          alt_vip_vfr_vga_avalon_streaming_source_ready;                         // alt_vip_itc_0:is_ready -> alt_vip_vfr_vga:dout_ready
	wire          alt_vip_vfr_vga_avalon_streaming_source_startofpacket;                 // alt_vip_vfr_vga:dout_startofpacket -> alt_vip_itc_0:is_sop
	wire          alt_vip_vfr_vga_avalon_streaming_source_endofpacket;                   // alt_vip_vfr_vga:dout_endofpacket -> alt_vip_itc_0:is_eop
	wire          fifo_dummy64_in_out_valid;                                             // fifo_dummy64_in:avalonst_source_valid -> fifo_dummy64_out:avalonst_sink_valid
	wire   [31:0] fifo_dummy64_in_out_data;                                              // fifo_dummy64_in:avalonst_source_data -> fifo_dummy64_out:avalonst_sink_data
	wire          fifo_dummy64_in_out_ready;                                             // fifo_dummy64_out:avalonst_sink_ready -> fifo_dummy64_in:avalonst_source_ready
	wire          gp_pll_outclk0_clk;                                                    // gp_pll:outclk_0 -> [alt_vip_itc_0:is_clk, alt_vip_vfr_vga:clock, mm_interconnect_1:gp_pll_outclk0_clk, rst_controller_002:clk]
	wire   [63:0] nmr_sys_pll_reconfig_from_pll_reconfig_from_pll;                       // nmr_sys_pll:reconfig_from_pll -> nmr_sys_pll_reconfig:reconfig_from_pll
	wire   [63:0] analyzer_pll_reconfig_from_pll_reconfig_from_pll;                      // analyzer_pll:reconfig_from_pll -> analyzer_pll_reconfig:reconfig_from_pll
	wire   [63:0] nmr_sys_pll_reconfig_reconfig_to_pll_reconfig_to_pll;                  // nmr_sys_pll_reconfig:reconfig_to_pll -> nmr_sys_pll:reconfig_to_pll
	wire   [63:0] analyzer_pll_reconfig_reconfig_to_pll_reconfig_to_pll;                 // analyzer_pll_reconfig:reconfig_to_pll -> analyzer_pll:reconfig_to_pll
	wire  [127:0] alt_vip_vfr_vga_avalon_master_readdata;                                // mm_interconnect_0:alt_vip_vfr_vga_avalon_master_readdata -> alt_vip_vfr_vga:master_readdata
	wire          alt_vip_vfr_vga_avalon_master_waitrequest;                             // mm_interconnect_0:alt_vip_vfr_vga_avalon_master_waitrequest -> alt_vip_vfr_vga:master_waitrequest
	wire   [31:0] alt_vip_vfr_vga_avalon_master_address;                                 // alt_vip_vfr_vga:master_address -> mm_interconnect_0:alt_vip_vfr_vga_avalon_master_address
	wire          alt_vip_vfr_vga_avalon_master_read;                                    // alt_vip_vfr_vga:master_read -> mm_interconnect_0:alt_vip_vfr_vga_avalon_master_read
	wire          alt_vip_vfr_vga_avalon_master_readdatavalid;                           // mm_interconnect_0:alt_vip_vfr_vga_avalon_master_readdatavalid -> alt_vip_vfr_vga:master_readdatavalid
	wire    [5:0] alt_vip_vfr_vga_avalon_master_burstcount;                              // alt_vip_vfr_vga:master_burstcount -> mm_interconnect_0:alt_vip_vfr_vga_avalon_master_burstcount
	wire   [31:0] master_secure_master_readdata;                                         // mm_interconnect_0:master_secure_master_readdata -> master_secure:master_readdata
	wire          master_secure_master_waitrequest;                                      // mm_interconnect_0:master_secure_master_waitrequest -> master_secure:master_waitrequest
	wire   [31:0] master_secure_master_address;                                          // master_secure:master_address -> mm_interconnect_0:master_secure_master_address
	wire          master_secure_master_read;                                             // master_secure:master_read -> mm_interconnect_0:master_secure_master_read
	wire    [3:0] master_secure_master_byteenable;                                       // master_secure:master_byteenable -> mm_interconnect_0:master_secure_master_byteenable
	wire          master_secure_master_readdatavalid;                                    // mm_interconnect_0:master_secure_master_readdatavalid -> master_secure:master_readdatavalid
	wire          master_secure_master_write;                                            // master_secure:master_write -> mm_interconnect_0:master_secure_master_write
	wire   [31:0] master_secure_master_writedata;                                        // master_secure:master_writedata -> mm_interconnect_0:master_secure_master_writedata
	wire    [1:0] mm_interconnect_0_hps_0_f2h_axi_slave_awburst;                         // mm_interconnect_0:hps_0_f2h_axi_slave_awburst -> hps_0:f2h_AWBURST
	wire    [4:0] mm_interconnect_0_hps_0_f2h_axi_slave_awuser;                          // mm_interconnect_0:hps_0_f2h_axi_slave_awuser -> hps_0:f2h_AWUSER
	wire    [3:0] mm_interconnect_0_hps_0_f2h_axi_slave_arlen;                           // mm_interconnect_0:hps_0_f2h_axi_slave_arlen -> hps_0:f2h_ARLEN
	wire   [15:0] mm_interconnect_0_hps_0_f2h_axi_slave_wstrb;                           // mm_interconnect_0:hps_0_f2h_axi_slave_wstrb -> hps_0:f2h_WSTRB
	wire          mm_interconnect_0_hps_0_f2h_axi_slave_wready;                          // hps_0:f2h_WREADY -> mm_interconnect_0:hps_0_f2h_axi_slave_wready
	wire    [7:0] mm_interconnect_0_hps_0_f2h_axi_slave_rid;                             // hps_0:f2h_RID -> mm_interconnect_0:hps_0_f2h_axi_slave_rid
	wire          mm_interconnect_0_hps_0_f2h_axi_slave_rready;                          // mm_interconnect_0:hps_0_f2h_axi_slave_rready -> hps_0:f2h_RREADY
	wire    [3:0] mm_interconnect_0_hps_0_f2h_axi_slave_awlen;                           // mm_interconnect_0:hps_0_f2h_axi_slave_awlen -> hps_0:f2h_AWLEN
	wire    [7:0] mm_interconnect_0_hps_0_f2h_axi_slave_wid;                             // mm_interconnect_0:hps_0_f2h_axi_slave_wid -> hps_0:f2h_WID
	wire    [3:0] mm_interconnect_0_hps_0_f2h_axi_slave_arcache;                         // mm_interconnect_0:hps_0_f2h_axi_slave_arcache -> hps_0:f2h_ARCACHE
	wire          mm_interconnect_0_hps_0_f2h_axi_slave_wvalid;                          // mm_interconnect_0:hps_0_f2h_axi_slave_wvalid -> hps_0:f2h_WVALID
	wire   [31:0] mm_interconnect_0_hps_0_f2h_axi_slave_araddr;                          // mm_interconnect_0:hps_0_f2h_axi_slave_araddr -> hps_0:f2h_ARADDR
	wire    [2:0] mm_interconnect_0_hps_0_f2h_axi_slave_arprot;                          // mm_interconnect_0:hps_0_f2h_axi_slave_arprot -> hps_0:f2h_ARPROT
	wire    [2:0] mm_interconnect_0_hps_0_f2h_axi_slave_awprot;                          // mm_interconnect_0:hps_0_f2h_axi_slave_awprot -> hps_0:f2h_AWPROT
	wire  [127:0] mm_interconnect_0_hps_0_f2h_axi_slave_wdata;                           // mm_interconnect_0:hps_0_f2h_axi_slave_wdata -> hps_0:f2h_WDATA
	wire          mm_interconnect_0_hps_0_f2h_axi_slave_arvalid;                         // mm_interconnect_0:hps_0_f2h_axi_slave_arvalid -> hps_0:f2h_ARVALID
	wire    [3:0] mm_interconnect_0_hps_0_f2h_axi_slave_awcache;                         // mm_interconnect_0:hps_0_f2h_axi_slave_awcache -> hps_0:f2h_AWCACHE
	wire    [7:0] mm_interconnect_0_hps_0_f2h_axi_slave_arid;                            // mm_interconnect_0:hps_0_f2h_axi_slave_arid -> hps_0:f2h_ARID
	wire    [1:0] mm_interconnect_0_hps_0_f2h_axi_slave_arlock;                          // mm_interconnect_0:hps_0_f2h_axi_slave_arlock -> hps_0:f2h_ARLOCK
	wire    [1:0] mm_interconnect_0_hps_0_f2h_axi_slave_awlock;                          // mm_interconnect_0:hps_0_f2h_axi_slave_awlock -> hps_0:f2h_AWLOCK
	wire   [31:0] mm_interconnect_0_hps_0_f2h_axi_slave_awaddr;                          // mm_interconnect_0:hps_0_f2h_axi_slave_awaddr -> hps_0:f2h_AWADDR
	wire    [1:0] mm_interconnect_0_hps_0_f2h_axi_slave_bresp;                           // hps_0:f2h_BRESP -> mm_interconnect_0:hps_0_f2h_axi_slave_bresp
	wire          mm_interconnect_0_hps_0_f2h_axi_slave_arready;                         // hps_0:f2h_ARREADY -> mm_interconnect_0:hps_0_f2h_axi_slave_arready
	wire  [127:0] mm_interconnect_0_hps_0_f2h_axi_slave_rdata;                           // hps_0:f2h_RDATA -> mm_interconnect_0:hps_0_f2h_axi_slave_rdata
	wire          mm_interconnect_0_hps_0_f2h_axi_slave_awready;                         // hps_0:f2h_AWREADY -> mm_interconnect_0:hps_0_f2h_axi_slave_awready
	wire    [1:0] mm_interconnect_0_hps_0_f2h_axi_slave_arburst;                         // mm_interconnect_0:hps_0_f2h_axi_slave_arburst -> hps_0:f2h_ARBURST
	wire    [2:0] mm_interconnect_0_hps_0_f2h_axi_slave_arsize;                          // mm_interconnect_0:hps_0_f2h_axi_slave_arsize -> hps_0:f2h_ARSIZE
	wire          mm_interconnect_0_hps_0_f2h_axi_slave_bready;                          // mm_interconnect_0:hps_0_f2h_axi_slave_bready -> hps_0:f2h_BREADY
	wire          mm_interconnect_0_hps_0_f2h_axi_slave_rlast;                           // hps_0:f2h_RLAST -> mm_interconnect_0:hps_0_f2h_axi_slave_rlast
	wire          mm_interconnect_0_hps_0_f2h_axi_slave_wlast;                           // mm_interconnect_0:hps_0_f2h_axi_slave_wlast -> hps_0:f2h_WLAST
	wire    [1:0] mm_interconnect_0_hps_0_f2h_axi_slave_rresp;                           // hps_0:f2h_RRESP -> mm_interconnect_0:hps_0_f2h_axi_slave_rresp
	wire    [7:0] mm_interconnect_0_hps_0_f2h_axi_slave_awid;                            // mm_interconnect_0:hps_0_f2h_axi_slave_awid -> hps_0:f2h_AWID
	wire    [7:0] mm_interconnect_0_hps_0_f2h_axi_slave_bid;                             // hps_0:f2h_BID -> mm_interconnect_0:hps_0_f2h_axi_slave_bid
	wire          mm_interconnect_0_hps_0_f2h_axi_slave_bvalid;                          // hps_0:f2h_BVALID -> mm_interconnect_0:hps_0_f2h_axi_slave_bvalid
	wire    [2:0] mm_interconnect_0_hps_0_f2h_axi_slave_awsize;                          // mm_interconnect_0:hps_0_f2h_axi_slave_awsize -> hps_0:f2h_AWSIZE
	wire          mm_interconnect_0_hps_0_f2h_axi_slave_awvalid;                         // mm_interconnect_0:hps_0_f2h_axi_slave_awvalid -> hps_0:f2h_AWVALID
	wire    [4:0] mm_interconnect_0_hps_0_f2h_axi_slave_aruser;                          // mm_interconnect_0:hps_0_f2h_axi_slave_aruser -> hps_0:f2h_ARUSER
	wire          mm_interconnect_0_hps_0_f2h_axi_slave_rvalid;                          // hps_0:f2h_RVALID -> mm_interconnect_0:hps_0_f2h_axi_slave_rvalid
	wire    [1:0] hps_0_h2f_axi_master_awburst;                                          // hps_0:h2f_AWBURST -> mm_interconnect_1:hps_0_h2f_axi_master_awburst
	wire    [3:0] hps_0_h2f_axi_master_arlen;                                            // hps_0:h2f_ARLEN -> mm_interconnect_1:hps_0_h2f_axi_master_arlen
	wire   [15:0] hps_0_h2f_axi_master_wstrb;                                            // hps_0:h2f_WSTRB -> mm_interconnect_1:hps_0_h2f_axi_master_wstrb
	wire          hps_0_h2f_axi_master_wready;                                           // mm_interconnect_1:hps_0_h2f_axi_master_wready -> hps_0:h2f_WREADY
	wire   [11:0] hps_0_h2f_axi_master_rid;                                              // mm_interconnect_1:hps_0_h2f_axi_master_rid -> hps_0:h2f_RID
	wire          hps_0_h2f_axi_master_rready;                                           // hps_0:h2f_RREADY -> mm_interconnect_1:hps_0_h2f_axi_master_rready
	wire    [3:0] hps_0_h2f_axi_master_awlen;                                            // hps_0:h2f_AWLEN -> mm_interconnect_1:hps_0_h2f_axi_master_awlen
	wire   [11:0] hps_0_h2f_axi_master_wid;                                              // hps_0:h2f_WID -> mm_interconnect_1:hps_0_h2f_axi_master_wid
	wire    [3:0] hps_0_h2f_axi_master_arcache;                                          // hps_0:h2f_ARCACHE -> mm_interconnect_1:hps_0_h2f_axi_master_arcache
	wire          hps_0_h2f_axi_master_wvalid;                                           // hps_0:h2f_WVALID -> mm_interconnect_1:hps_0_h2f_axi_master_wvalid
	wire   [29:0] hps_0_h2f_axi_master_araddr;                                           // hps_0:h2f_ARADDR -> mm_interconnect_1:hps_0_h2f_axi_master_araddr
	wire    [2:0] hps_0_h2f_axi_master_arprot;                                           // hps_0:h2f_ARPROT -> mm_interconnect_1:hps_0_h2f_axi_master_arprot
	wire    [2:0] hps_0_h2f_axi_master_awprot;                                           // hps_0:h2f_AWPROT -> mm_interconnect_1:hps_0_h2f_axi_master_awprot
	wire  [127:0] hps_0_h2f_axi_master_wdata;                                            // hps_0:h2f_WDATA -> mm_interconnect_1:hps_0_h2f_axi_master_wdata
	wire          hps_0_h2f_axi_master_arvalid;                                          // hps_0:h2f_ARVALID -> mm_interconnect_1:hps_0_h2f_axi_master_arvalid
	wire    [3:0] hps_0_h2f_axi_master_awcache;                                          // hps_0:h2f_AWCACHE -> mm_interconnect_1:hps_0_h2f_axi_master_awcache
	wire   [11:0] hps_0_h2f_axi_master_arid;                                             // hps_0:h2f_ARID -> mm_interconnect_1:hps_0_h2f_axi_master_arid
	wire    [1:0] hps_0_h2f_axi_master_arlock;                                           // hps_0:h2f_ARLOCK -> mm_interconnect_1:hps_0_h2f_axi_master_arlock
	wire    [1:0] hps_0_h2f_axi_master_awlock;                                           // hps_0:h2f_AWLOCK -> mm_interconnect_1:hps_0_h2f_axi_master_awlock
	wire   [29:0] hps_0_h2f_axi_master_awaddr;                                           // hps_0:h2f_AWADDR -> mm_interconnect_1:hps_0_h2f_axi_master_awaddr
	wire    [1:0] hps_0_h2f_axi_master_bresp;                                            // mm_interconnect_1:hps_0_h2f_axi_master_bresp -> hps_0:h2f_BRESP
	wire          hps_0_h2f_axi_master_arready;                                          // mm_interconnect_1:hps_0_h2f_axi_master_arready -> hps_0:h2f_ARREADY
	wire  [127:0] hps_0_h2f_axi_master_rdata;                                            // mm_interconnect_1:hps_0_h2f_axi_master_rdata -> hps_0:h2f_RDATA
	wire          hps_0_h2f_axi_master_awready;                                          // mm_interconnect_1:hps_0_h2f_axi_master_awready -> hps_0:h2f_AWREADY
	wire    [1:0] hps_0_h2f_axi_master_arburst;                                          // hps_0:h2f_ARBURST -> mm_interconnect_1:hps_0_h2f_axi_master_arburst
	wire    [2:0] hps_0_h2f_axi_master_arsize;                                           // hps_0:h2f_ARSIZE -> mm_interconnect_1:hps_0_h2f_axi_master_arsize
	wire          hps_0_h2f_axi_master_bready;                                           // hps_0:h2f_BREADY -> mm_interconnect_1:hps_0_h2f_axi_master_bready
	wire          hps_0_h2f_axi_master_rlast;                                            // mm_interconnect_1:hps_0_h2f_axi_master_rlast -> hps_0:h2f_RLAST
	wire          hps_0_h2f_axi_master_wlast;                                            // hps_0:h2f_WLAST -> mm_interconnect_1:hps_0_h2f_axi_master_wlast
	wire    [1:0] hps_0_h2f_axi_master_rresp;                                            // mm_interconnect_1:hps_0_h2f_axi_master_rresp -> hps_0:h2f_RRESP
	wire   [11:0] hps_0_h2f_axi_master_awid;                                             // hps_0:h2f_AWID -> mm_interconnect_1:hps_0_h2f_axi_master_awid
	wire   [11:0] hps_0_h2f_axi_master_bid;                                              // mm_interconnect_1:hps_0_h2f_axi_master_bid -> hps_0:h2f_BID
	wire          hps_0_h2f_axi_master_bvalid;                                           // mm_interconnect_1:hps_0_h2f_axi_master_bvalid -> hps_0:h2f_BVALID
	wire    [2:0] hps_0_h2f_axi_master_awsize;                                           // hps_0:h2f_AWSIZE -> mm_interconnect_1:hps_0_h2f_axi_master_awsize
	wire          hps_0_h2f_axi_master_awvalid;                                          // hps_0:h2f_AWVALID -> mm_interconnect_1:hps_0_h2f_axi_master_awvalid
	wire          hps_0_h2f_axi_master_rvalid;                                           // mm_interconnect_1:hps_0_h2f_axi_master_rvalid -> hps_0:h2f_RVALID
	wire          dma_fifo_write_master_chipselect;                                      // dma_fifo:write_chipselect -> mm_interconnect_1:dma_fifo_write_master_chipselect
	wire          dma_fifo_write_master_waitrequest;                                     // mm_interconnect_1:dma_fifo_write_master_waitrequest -> dma_fifo:write_waitrequest
	wire   [25:0] dma_fifo_write_master_address;                                         // dma_fifo:write_address -> mm_interconnect_1:dma_fifo_write_master_address
	wire    [3:0] dma_fifo_write_master_byteenable;                                      // dma_fifo:write_byteenable -> mm_interconnect_1:dma_fifo_write_master_byteenable
	wire          dma_fifo_write_master_write;                                           // dma_fifo:write_write_n -> mm_interconnect_1:dma_fifo_write_master_write
	wire   [31:0] dma_fifo_write_master_writedata;                                       // dma_fifo:write_writedata -> mm_interconnect_1:dma_fifo_write_master_writedata
	wire          dma_dconvi_write_master_chipselect;                                    // dma_dconvi:write_chipselect -> mm_interconnect_1:dma_dconvi_write_master_chipselect
	wire          dma_dconvi_write_master_waitrequest;                                   // mm_interconnect_1:dma_dconvi_write_master_waitrequest -> dma_dconvi:write_waitrequest
	wire   [25:0] dma_dconvi_write_master_address;                                       // dma_dconvi:write_address -> mm_interconnect_1:dma_dconvi_write_master_address
	wire    [3:0] dma_dconvi_write_master_byteenable;                                    // dma_dconvi:write_byteenable -> mm_interconnect_1:dma_dconvi_write_master_byteenable
	wire          dma_dconvi_write_master_write;                                         // dma_dconvi:write_write_n -> mm_interconnect_1:dma_dconvi_write_master_write
	wire   [31:0] dma_dconvi_write_master_writedata;                                     // dma_dconvi:write_writedata -> mm_interconnect_1:dma_dconvi_write_master_writedata
	wire          dma_dconvq_write_master_chipselect;                                    // dma_dconvq:write_chipselect -> mm_interconnect_1:dma_dconvq_write_master_chipselect
	wire          dma_dconvq_write_master_waitrequest;                                   // mm_interconnect_1:dma_dconvq_write_master_waitrequest -> dma_dconvq:write_waitrequest
	wire   [25:0] dma_dconvq_write_master_address;                                       // dma_dconvq:write_address -> mm_interconnect_1:dma_dconvq_write_master_address
	wire    [3:0] dma_dconvq_write_master_byteenable;                                    // dma_dconvq:write_byteenable -> mm_interconnect_1:dma_dconvq_write_master_byteenable
	wire          dma_dconvq_write_master_write;                                         // dma_dconvq:write_write_n -> mm_interconnect_1:dma_dconvq_write_master_write
	wire   [31:0] dma_dconvq_write_master_writedata;                                     // dma_dconvq:write_writedata -> mm_interconnect_1:dma_dconvq_write_master_writedata
	wire          dma_dummy_write_master_chipselect;                                     // dma_dummy:write_chipselect -> mm_interconnect_1:dma_dummy_write_master_chipselect
	wire          dma_dummy_write_master_waitrequest;                                    // mm_interconnect_1:dma_dummy_write_master_waitrequest -> dma_dummy:write_waitrequest
	wire   [25:0] dma_dummy_write_master_address;                                        // dma_dummy:write_address -> mm_interconnect_1:dma_dummy_write_master_address
	wire    [3:0] dma_dummy_write_master_byteenable;                                     // dma_dummy:write_byteenable -> mm_interconnect_1:dma_dummy_write_master_byteenable
	wire          dma_dummy_write_master_write;                                          // dma_dummy:write_write_n -> mm_interconnect_1:dma_dummy_write_master_write
	wire   [31:0] dma_dummy_write_master_writedata;                                      // dma_dummy:write_writedata -> mm_interconnect_1:dma_dummy_write_master_writedata
	wire          dma_fifo_read_master_chipselect;                                       // dma_fifo:read_chipselect -> mm_interconnect_1:dma_fifo_read_master_chipselect
	wire   [31:0] dma_fifo_read_master_readdata;                                         // mm_interconnect_1:dma_fifo_read_master_readdata -> dma_fifo:read_readdata
	wire          dma_fifo_read_master_waitrequest;                                      // mm_interconnect_1:dma_fifo_read_master_waitrequest -> dma_fifo:read_waitrequest
	wire   [26:0] dma_fifo_read_master_address;                                          // dma_fifo:read_address -> mm_interconnect_1:dma_fifo_read_master_address
	wire          dma_fifo_read_master_read;                                             // dma_fifo:read_read_n -> mm_interconnect_1:dma_fifo_read_master_read
	wire          dma_fifo_read_master_readdatavalid;                                    // mm_interconnect_1:dma_fifo_read_master_readdatavalid -> dma_fifo:read_readdatavalid
	wire    [1:0] hps_0_h2f_lw_axi_master_awburst;                                       // hps_0:h2f_lw_AWBURST -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awburst
	wire    [3:0] hps_0_h2f_lw_axi_master_arlen;                                         // hps_0:h2f_lw_ARLEN -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arlen
	wire    [3:0] hps_0_h2f_lw_axi_master_wstrb;                                         // hps_0:h2f_lw_WSTRB -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wstrb
	wire          hps_0_h2f_lw_axi_master_wready;                                        // mm_interconnect_1:hps_0_h2f_lw_axi_master_wready -> hps_0:h2f_lw_WREADY
	wire   [11:0] hps_0_h2f_lw_axi_master_rid;                                           // mm_interconnect_1:hps_0_h2f_lw_axi_master_rid -> hps_0:h2f_lw_RID
	wire          hps_0_h2f_lw_axi_master_rready;                                        // hps_0:h2f_lw_RREADY -> mm_interconnect_1:hps_0_h2f_lw_axi_master_rready
	wire    [3:0] hps_0_h2f_lw_axi_master_awlen;                                         // hps_0:h2f_lw_AWLEN -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awlen
	wire   [11:0] hps_0_h2f_lw_axi_master_wid;                                           // hps_0:h2f_lw_WID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wid
	wire    [3:0] hps_0_h2f_lw_axi_master_arcache;                                       // hps_0:h2f_lw_ARCACHE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arcache
	wire          hps_0_h2f_lw_axi_master_wvalid;                                        // hps_0:h2f_lw_WVALID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wvalid
	wire   [20:0] hps_0_h2f_lw_axi_master_araddr;                                        // hps_0:h2f_lw_ARADDR -> mm_interconnect_1:hps_0_h2f_lw_axi_master_araddr
	wire    [2:0] hps_0_h2f_lw_axi_master_arprot;                                        // hps_0:h2f_lw_ARPROT -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arprot
	wire    [2:0] hps_0_h2f_lw_axi_master_awprot;                                        // hps_0:h2f_lw_AWPROT -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awprot
	wire   [31:0] hps_0_h2f_lw_axi_master_wdata;                                         // hps_0:h2f_lw_WDATA -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wdata
	wire          hps_0_h2f_lw_axi_master_arvalid;                                       // hps_0:h2f_lw_ARVALID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arvalid
	wire    [3:0] hps_0_h2f_lw_axi_master_awcache;                                       // hps_0:h2f_lw_AWCACHE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awcache
	wire   [11:0] hps_0_h2f_lw_axi_master_arid;                                          // hps_0:h2f_lw_ARID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arid
	wire    [1:0] hps_0_h2f_lw_axi_master_arlock;                                        // hps_0:h2f_lw_ARLOCK -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arlock
	wire    [1:0] hps_0_h2f_lw_axi_master_awlock;                                        // hps_0:h2f_lw_AWLOCK -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awlock
	wire   [20:0] hps_0_h2f_lw_axi_master_awaddr;                                        // hps_0:h2f_lw_AWADDR -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awaddr
	wire    [1:0] hps_0_h2f_lw_axi_master_bresp;                                         // mm_interconnect_1:hps_0_h2f_lw_axi_master_bresp -> hps_0:h2f_lw_BRESP
	wire          hps_0_h2f_lw_axi_master_arready;                                       // mm_interconnect_1:hps_0_h2f_lw_axi_master_arready -> hps_0:h2f_lw_ARREADY
	wire   [31:0] hps_0_h2f_lw_axi_master_rdata;                                         // mm_interconnect_1:hps_0_h2f_lw_axi_master_rdata -> hps_0:h2f_lw_RDATA
	wire          hps_0_h2f_lw_axi_master_awready;                                       // mm_interconnect_1:hps_0_h2f_lw_axi_master_awready -> hps_0:h2f_lw_AWREADY
	wire    [1:0] hps_0_h2f_lw_axi_master_arburst;                                       // hps_0:h2f_lw_ARBURST -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arburst
	wire    [2:0] hps_0_h2f_lw_axi_master_arsize;                                        // hps_0:h2f_lw_ARSIZE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arsize
	wire          hps_0_h2f_lw_axi_master_bready;                                        // hps_0:h2f_lw_BREADY -> mm_interconnect_1:hps_0_h2f_lw_axi_master_bready
	wire          hps_0_h2f_lw_axi_master_rlast;                                         // mm_interconnect_1:hps_0_h2f_lw_axi_master_rlast -> hps_0:h2f_lw_RLAST
	wire          hps_0_h2f_lw_axi_master_wlast;                                         // hps_0:h2f_lw_WLAST -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wlast
	wire    [1:0] hps_0_h2f_lw_axi_master_rresp;                                         // mm_interconnect_1:hps_0_h2f_lw_axi_master_rresp -> hps_0:h2f_lw_RRESP
	wire   [11:0] hps_0_h2f_lw_axi_master_awid;                                          // hps_0:h2f_lw_AWID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awid
	wire   [11:0] hps_0_h2f_lw_axi_master_bid;                                           // mm_interconnect_1:hps_0_h2f_lw_axi_master_bid -> hps_0:h2f_lw_BID
	wire          hps_0_h2f_lw_axi_master_bvalid;                                        // mm_interconnect_1:hps_0_h2f_lw_axi_master_bvalid -> hps_0:h2f_lw_BVALID
	wire    [2:0] hps_0_h2f_lw_axi_master_awsize;                                        // hps_0:h2f_lw_AWSIZE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awsize
	wire          hps_0_h2f_lw_axi_master_awvalid;                                       // hps_0:h2f_lw_AWVALID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awvalid
	wire          hps_0_h2f_lw_axi_master_rvalid;                                        // mm_interconnect_1:hps_0_h2f_lw_axi_master_rvalid -> hps_0:h2f_lw_RVALID
	wire   [31:0] master_non_sec_master_readdata;                                        // mm_interconnect_1:master_non_sec_master_readdata -> master_non_sec:master_readdata
	wire          master_non_sec_master_waitrequest;                                     // mm_interconnect_1:master_non_sec_master_waitrequest -> master_non_sec:master_waitrequest
	wire   [31:0] master_non_sec_master_address;                                         // master_non_sec:master_address -> mm_interconnect_1:master_non_sec_master_address
	wire          master_non_sec_master_read;                                            // master_non_sec:master_read -> mm_interconnect_1:master_non_sec_master_read
	wire    [3:0] master_non_sec_master_byteenable;                                      // master_non_sec:master_byteenable -> mm_interconnect_1:master_non_sec_master_byteenable
	wire          master_non_sec_master_readdatavalid;                                   // mm_interconnect_1:master_non_sec_master_readdatavalid -> master_non_sec:master_readdatavalid
	wire          master_non_sec_master_write;                                           // master_non_sec:master_write -> mm_interconnect_1:master_non_sec_master_write
	wire   [31:0] master_non_sec_master_writedata;                                       // master_non_sec:master_writedata -> mm_interconnect_1:master_non_sec_master_writedata
	wire          dma_dconvq_read_master_chipselect;                                     // dma_dconvq:read_chipselect -> mm_interconnect_1:dma_dconvq_read_master_chipselect
	wire   [31:0] dma_dconvq_read_master_readdata;                                       // mm_interconnect_1:dma_dconvq_read_master_readdata -> dma_dconvq:read_readdata
	wire          dma_dconvq_read_master_waitrequest;                                    // mm_interconnect_1:dma_dconvq_read_master_waitrequest -> dma_dconvq:read_waitrequest
	wire   [10:0] dma_dconvq_read_master_address;                                        // dma_dconvq:read_address -> mm_interconnect_1:dma_dconvq_read_master_address
	wire          dma_dconvq_read_master_read;                                           // dma_dconvq:read_read_n -> mm_interconnect_1:dma_dconvq_read_master_read
	wire          dma_dconvq_read_master_readdatavalid;                                  // mm_interconnect_1:dma_dconvq_read_master_readdatavalid -> dma_dconvq:read_readdatavalid
	wire          dma_dconvi_read_master_chipselect;                                     // dma_dconvi:read_chipselect -> mm_interconnect_1:dma_dconvi_read_master_chipselect
	wire   [31:0] dma_dconvi_read_master_readdata;                                       // mm_interconnect_1:dma_dconvi_read_master_readdata -> dma_dconvi:read_readdata
	wire          dma_dconvi_read_master_waitrequest;                                    // mm_interconnect_1:dma_dconvi_read_master_waitrequest -> dma_dconvi:read_waitrequest
	wire   [10:0] dma_dconvi_read_master_address;                                        // dma_dconvi:read_address -> mm_interconnect_1:dma_dconvi_read_master_address
	wire          dma_dconvi_read_master_read;                                           // dma_dconvi:read_read_n -> mm_interconnect_1:dma_dconvi_read_master_read
	wire          dma_dconvi_read_master_readdatavalid;                                  // mm_interconnect_1:dma_dconvi_read_master_readdatavalid -> dma_dconvi:read_readdatavalid
	wire          dma_dummy_read_master_chipselect;                                      // dma_dummy:read_chipselect -> mm_interconnect_1:dma_dummy_read_master_chipselect
	wire   [31:0] dma_dummy_read_master_readdata;                                        // mm_interconnect_1:dma_dummy_read_master_readdata -> dma_dummy:read_readdata
	wire          dma_dummy_read_master_waitrequest;                                     // mm_interconnect_1:dma_dummy_read_master_waitrequest -> dma_dummy:read_waitrequest
	wire   [26:0] dma_dummy_read_master_address;                                         // dma_dummy:read_address -> mm_interconnect_1:dma_dummy_read_master_address
	wire          dma_dummy_read_master_read;                                            // dma_dummy:read_read_n -> mm_interconnect_1:dma_dummy_read_master_read
	wire          dma_dummy_read_master_readdatavalid;                                   // mm_interconnect_1:dma_dummy_read_master_readdatavalid -> dma_dummy:read_readdatavalid
	wire          mm_interconnect_1_fifo_dummy64_in_in_waitrequest;                      // fifo_dummy64_in:avalonmm_write_slave_waitrequest -> mm_interconnect_1:fifo_dummy64_in_in_waitrequest
	wire    [0:0] mm_interconnect_1_fifo_dummy64_in_in_address;                          // mm_interconnect_1:fifo_dummy64_in_in_address -> fifo_dummy64_in:avalonmm_write_slave_address
	wire          mm_interconnect_1_fifo_dummy64_in_in_write;                            // mm_interconnect_1:fifo_dummy64_in_in_write -> fifo_dummy64_in:avalonmm_write_slave_write
	wire   [31:0] mm_interconnect_1_fifo_dummy64_in_in_writedata;                        // mm_interconnect_1:fifo_dummy64_in_in_writedata -> fifo_dummy64_in:avalonmm_write_slave_writedata
	wire          mm_interconnect_1_fifo_dummy_in_waitrequest;                           // fifo_dummy:avalonmm_write_slave_waitrequest -> mm_interconnect_1:fifo_dummy_in_waitrequest
	wire          mm_interconnect_1_fifo_dummy_in_write;                                 // mm_interconnect_1:fifo_dummy_in_write -> fifo_dummy:avalonmm_write_slave_write
	wire   [31:0] mm_interconnect_1_fifo_dummy_in_writedata;                             // mm_interconnect_1:fifo_dummy_in_writedata -> fifo_dummy:avalonmm_write_slave_writedata
	wire   [31:0] mm_interconnect_1_fifo_dummy64_in_in_csr_readdata;                     // fifo_dummy64_in:wrclk_control_slave_readdata -> mm_interconnect_1:fifo_dummy64_in_in_csr_readdata
	wire    [2:0] mm_interconnect_1_fifo_dummy64_in_in_csr_address;                      // mm_interconnect_1:fifo_dummy64_in_in_csr_address -> fifo_dummy64_in:wrclk_control_slave_address
	wire          mm_interconnect_1_fifo_dummy64_in_in_csr_read;                         // mm_interconnect_1:fifo_dummy64_in_in_csr_read -> fifo_dummy64_in:wrclk_control_slave_read
	wire          mm_interconnect_1_fifo_dummy64_in_in_csr_write;                        // mm_interconnect_1:fifo_dummy64_in_in_csr_write -> fifo_dummy64_in:wrclk_control_slave_write
	wire   [31:0] mm_interconnect_1_fifo_dummy64_in_in_csr_writedata;                    // mm_interconnect_1:fifo_dummy64_in_in_csr_writedata -> fifo_dummy64_in:wrclk_control_slave_writedata
	wire   [31:0] mm_interconnect_1_fifo_dummy64_out_in_csr_readdata;                    // fifo_dummy64_out:wrclk_control_slave_readdata -> mm_interconnect_1:fifo_dummy64_out_in_csr_readdata
	wire    [2:0] mm_interconnect_1_fifo_dummy64_out_in_csr_address;                     // mm_interconnect_1:fifo_dummy64_out_in_csr_address -> fifo_dummy64_out:wrclk_control_slave_address
	wire          mm_interconnect_1_fifo_dummy64_out_in_csr_read;                        // mm_interconnect_1:fifo_dummy64_out_in_csr_read -> fifo_dummy64_out:wrclk_control_slave_read
	wire          mm_interconnect_1_fifo_dummy64_out_in_csr_write;                       // mm_interconnect_1:fifo_dummy64_out_in_csr_write -> fifo_dummy64_out:wrclk_control_slave_write
	wire   [31:0] mm_interconnect_1_fifo_dummy64_out_in_csr_writedata;                   // mm_interconnect_1:fifo_dummy64_out_in_csr_writedata -> fifo_dummy64_out:wrclk_control_slave_writedata
	wire   [31:0] mm_interconnect_1_fifo_dummy_in_csr_readdata;                          // fifo_dummy:wrclk_control_slave_readdata -> mm_interconnect_1:fifo_dummy_in_csr_readdata
	wire    [2:0] mm_interconnect_1_fifo_dummy_in_csr_address;                           // mm_interconnect_1:fifo_dummy_in_csr_address -> fifo_dummy:wrclk_control_slave_address
	wire          mm_interconnect_1_fifo_dummy_in_csr_read;                              // mm_interconnect_1:fifo_dummy_in_csr_read -> fifo_dummy:wrclk_control_slave_read
	wire          mm_interconnect_1_fifo_dummy_in_csr_write;                             // mm_interconnect_1:fifo_dummy_in_csr_write -> fifo_dummy:wrclk_control_slave_write
	wire   [31:0] mm_interconnect_1_fifo_dummy_in_csr_writedata;                         // mm_interconnect_1:fifo_dummy_in_csr_writedata -> fifo_dummy:wrclk_control_slave_writedata
	wire   [31:0] mm_interconnect_1_fifo_dummy64_out_out_readdata;                       // fifo_dummy64_out:avalonmm_read_slave_readdata -> mm_interconnect_1:fifo_dummy64_out_out_readdata
	wire          mm_interconnect_1_fifo_dummy64_out_out_waitrequest;                    // fifo_dummy64_out:avalonmm_read_slave_waitrequest -> mm_interconnect_1:fifo_dummy64_out_out_waitrequest
	wire    [0:0] mm_interconnect_1_fifo_dummy64_out_out_address;                        // mm_interconnect_1:fifo_dummy64_out_out_address -> fifo_dummy64_out:avalonmm_read_slave_address
	wire          mm_interconnect_1_fifo_dummy64_out_out_read;                           // mm_interconnect_1:fifo_dummy64_out_out_read -> fifo_dummy64_out:avalonmm_read_slave_read
	wire   [31:0] mm_interconnect_1_fifo_dummy_out_readdata;                             // fifo_dummy:avalonmm_read_slave_readdata -> mm_interconnect_1:fifo_dummy_out_readdata
	wire          mm_interconnect_1_fifo_dummy_out_waitrequest;                          // fifo_dummy:avalonmm_read_slave_waitrequest -> mm_interconnect_1:fifo_dummy_out_waitrequest
	wire          mm_interconnect_1_fifo_dummy_out_read;                                 // mm_interconnect_1:fifo_dummy_out_read -> fifo_dummy:avalonmm_read_slave_read
	wire   [31:0] mm_interconnect_1_switches_s1_readdata;                                // switches:readdata -> mm_interconnect_1:switches_s1_readdata
	wire    [1:0] mm_interconnect_1_switches_s1_address;                                 // mm_interconnect_1:switches_s1_address -> switches:address
	wire          mm_interconnect_1_sdram_s1_chipselect;                                 // mm_interconnect_1:sdram_s1_chipselect -> sdram:az_cs
	wire   [15:0] mm_interconnect_1_sdram_s1_readdata;                                   // sdram:za_data -> mm_interconnect_1:sdram_s1_readdata
	wire          mm_interconnect_1_sdram_s1_waitrequest;                                // sdram:za_waitrequest -> mm_interconnect_1:sdram_s1_waitrequest
	wire   [24:0] mm_interconnect_1_sdram_s1_address;                                    // mm_interconnect_1:sdram_s1_address -> sdram:az_addr
	wire          mm_interconnect_1_sdram_s1_read;                                       // mm_interconnect_1:sdram_s1_read -> sdram:az_rd_n
	wire    [1:0] mm_interconnect_1_sdram_s1_byteenable;                                 // mm_interconnect_1:sdram_s1_byteenable -> sdram:az_be_n
	wire          mm_interconnect_1_sdram_s1_readdatavalid;                              // sdram:za_valid -> mm_interconnect_1:sdram_s1_readdatavalid
	wire          mm_interconnect_1_sdram_s1_write;                                      // mm_interconnect_1:sdram_s1_write -> sdram:az_wr_n
	wire   [15:0] mm_interconnect_1_sdram_s1_writedata;                                  // mm_interconnect_1:sdram_s1_writedata -> sdram:az_data
	wire   [31:0] mm_interconnect_1_adc_fifo_mem_out_readdata;                           // adc_fifo_mem:avalonmm_read_slave_readdata -> mm_interconnect_1:adc_fifo_mem_out_readdata
	wire          mm_interconnect_1_adc_fifo_mem_out_waitrequest;                        // adc_fifo_mem:avalonmm_read_slave_waitrequest -> mm_interconnect_1:adc_fifo_mem_out_waitrequest
	wire    [0:0] mm_interconnect_1_adc_fifo_mem_out_address;                            // mm_interconnect_1:adc_fifo_mem_out_address -> adc_fifo_mem:avalonmm_read_slave_address
	wire          mm_interconnect_1_adc_fifo_mem_out_read;                               // mm_interconnect_1:adc_fifo_mem_out_read -> adc_fifo_mem:avalonmm_read_slave_read
	wire          mm_interconnect_1_nmr_parameters_adc_val_sub_s1_chipselect;            // mm_interconnect_1:nmr_parameters_adc_val_sub_s1_chipselect -> nmr_parameters:adc_val_sub_s1_chipselect
	wire   [31:0] mm_interconnect_1_nmr_parameters_adc_val_sub_s1_readdata;              // nmr_parameters:adc_val_sub_s1_readdata -> mm_interconnect_1:nmr_parameters_adc_val_sub_s1_readdata
	wire    [1:0] mm_interconnect_1_nmr_parameters_adc_val_sub_s1_address;               // mm_interconnect_1:nmr_parameters_adc_val_sub_s1_address -> nmr_parameters:adc_val_sub_s1_address
	wire          mm_interconnect_1_nmr_parameters_adc_val_sub_s1_write;                 // mm_interconnect_1:nmr_parameters_adc_val_sub_s1_write -> nmr_parameters:adc_val_sub_s1_write_n
	wire   [31:0] mm_interconnect_1_nmr_parameters_adc_val_sub_s1_writedata;             // mm_interconnect_1:nmr_parameters_adc_val_sub_s1_writedata -> nmr_parameters:adc_val_sub_s1_writedata
	wire          mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect;              // mm_interconnect_1:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire   [31:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata;                // jtag_uart:av_readdata -> mm_interconnect_1:jtag_uart_avalon_jtag_slave_readdata
	wire          mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest;             // jtag_uart:av_waitrequest -> mm_interconnect_1:jtag_uart_avalon_jtag_slave_waitrequest
	wire    [0:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_address;                 // mm_interconnect_1:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire          mm_interconnect_1_jtag_uart_avalon_jtag_slave_read;                    // mm_interconnect_1:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire          mm_interconnect_1_jtag_uart_avalon_jtag_slave_write;                   // mm_interconnect_1:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire   [31:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata;               // mm_interconnect_1:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire   [15:0] mm_interconnect_1_dconv_fir_avalon_mm_slave_readdata;                  // dconv_fir:coeff_out_data -> mm_interconnect_1:dconv_fir_avalon_mm_slave_readdata
	wire    [5:0] mm_interconnect_1_dconv_fir_avalon_mm_slave_address;                   // mm_interconnect_1:dconv_fir_avalon_mm_slave_address -> dconv_fir:coeff_in_address
	wire          mm_interconnect_1_dconv_fir_avalon_mm_slave_read;                      // mm_interconnect_1:dconv_fir_avalon_mm_slave_read -> dconv_fir:coeff_in_read
	wire          mm_interconnect_1_dconv_fir_avalon_mm_slave_readdatavalid;             // dconv_fir:coeff_out_valid -> mm_interconnect_1:dconv_fir_avalon_mm_slave_readdatavalid
	wire          mm_interconnect_1_dconv_fir_avalon_mm_slave_write;                     // mm_interconnect_1:dconv_fir_avalon_mm_slave_write -> dconv_fir:coeff_in_we
	wire   [15:0] mm_interconnect_1_dconv_fir_avalon_mm_slave_writedata;                 // mm_interconnect_1:dconv_fir_avalon_mm_slave_writedata -> dconv_fir:coeff_in_data
	wire   [15:0] mm_interconnect_1_dconv_fir_q_avalon_mm_slave_readdata;                // dconv_fir_q:coeff_out_data -> mm_interconnect_1:dconv_fir_q_avalon_mm_slave_readdata
	wire    [5:0] mm_interconnect_1_dconv_fir_q_avalon_mm_slave_address;                 // mm_interconnect_1:dconv_fir_q_avalon_mm_slave_address -> dconv_fir_q:coeff_in_address
	wire          mm_interconnect_1_dconv_fir_q_avalon_mm_slave_read;                    // mm_interconnect_1:dconv_fir_q_avalon_mm_slave_read -> dconv_fir_q:coeff_in_read
	wire          mm_interconnect_1_dconv_fir_q_avalon_mm_slave_readdatavalid;           // dconv_fir_q:coeff_out_valid -> mm_interconnect_1:dconv_fir_q_avalon_mm_slave_readdatavalid
	wire          mm_interconnect_1_dconv_fir_q_avalon_mm_slave_write;                   // mm_interconnect_1:dconv_fir_q_avalon_mm_slave_write -> dconv_fir_q:coeff_in_we
	wire   [15:0] mm_interconnect_1_dconv_fir_q_avalon_mm_slave_writedata;               // mm_interconnect_1:dconv_fir_q_avalon_mm_slave_writedata -> dconv_fir_q:coeff_in_data
	wire   [31:0] mm_interconnect_1_alt_vip_vfr_vga_avalon_slave_readdata;               // alt_vip_vfr_vga:slave_readdata -> mm_interconnect_1:alt_vip_vfr_vga_avalon_slave_readdata
	wire    [4:0] mm_interconnect_1_alt_vip_vfr_vga_avalon_slave_address;                // mm_interconnect_1:alt_vip_vfr_vga_avalon_slave_address -> alt_vip_vfr_vga:slave_address
	wire          mm_interconnect_1_alt_vip_vfr_vga_avalon_slave_read;                   // mm_interconnect_1:alt_vip_vfr_vga_avalon_slave_read -> alt_vip_vfr_vga:slave_read
	wire          mm_interconnect_1_alt_vip_vfr_vga_avalon_slave_write;                  // mm_interconnect_1:alt_vip_vfr_vga_avalon_slave_write -> alt_vip_vfr_vga:slave_write
	wire   [31:0] mm_interconnect_1_alt_vip_vfr_vga_avalon_slave_writedata;              // mm_interconnect_1:alt_vip_vfr_vga_avalon_slave_writedata -> alt_vip_vfr_vga:slave_writedata
	wire   [31:0] mm_interconnect_1_sysid_qsys_control_slave_readdata;                   // sysid_qsys:readdata -> mm_interconnect_1:sysid_qsys_control_slave_readdata
	wire    [0:0] mm_interconnect_1_sysid_qsys_control_slave_address;                    // mm_interconnect_1:sysid_qsys_control_slave_address -> sysid_qsys:address
	wire   [31:0] mm_interconnect_1_i2c_int_csr_readdata;                                // i2c_int:readdata -> mm_interconnect_1:i2c_int_csr_readdata
	wire    [3:0] mm_interconnect_1_i2c_int_csr_address;                                 // mm_interconnect_1:i2c_int_csr_address -> i2c_int:addr
	wire          mm_interconnect_1_i2c_int_csr_read;                                    // mm_interconnect_1:i2c_int_csr_read -> i2c_int:read
	wire          mm_interconnect_1_i2c_int_csr_write;                                   // mm_interconnect_1:i2c_int_csr_write -> i2c_int:write
	wire   [31:0] mm_interconnect_1_i2c_int_csr_writedata;                               // mm_interconnect_1:i2c_int_csr_writedata -> i2c_int:writedata
	wire   [31:0] mm_interconnect_1_i2c_ext_csr_readdata;                                // i2c_ext:readdata -> mm_interconnect_1:i2c_ext_csr_readdata
	wire    [3:0] mm_interconnect_1_i2c_ext_csr_address;                                 // mm_interconnect_1:i2c_ext_csr_address -> i2c_ext:addr
	wire          mm_interconnect_1_i2c_ext_csr_read;                                    // mm_interconnect_1:i2c_ext_csr_read -> i2c_ext:read
	wire          mm_interconnect_1_i2c_ext_csr_write;                                   // mm_interconnect_1:i2c_ext_csr_write -> i2c_ext:write
	wire   [31:0] mm_interconnect_1_i2c_ext_csr_writedata;                               // mm_interconnect_1:i2c_ext_csr_writedata -> i2c_ext:writedata
	wire          mm_interconnect_1_nmr_parameters_delay_nosig_s1_chipselect;            // mm_interconnect_1:nmr_parameters_delay_nosig_s1_chipselect -> nmr_parameters:delay_nosig_s1_chipselect
	wire   [31:0] mm_interconnect_1_nmr_parameters_delay_nosig_s1_readdata;              // nmr_parameters:delay_nosig_s1_readdata -> mm_interconnect_1:nmr_parameters_delay_nosig_s1_readdata
	wire    [1:0] mm_interconnect_1_nmr_parameters_delay_nosig_s1_address;               // mm_interconnect_1:nmr_parameters_delay_nosig_s1_address -> nmr_parameters:delay_nosig_s1_address
	wire          mm_interconnect_1_nmr_parameters_delay_nosig_s1_write;                 // mm_interconnect_1:nmr_parameters_delay_nosig_s1_write -> nmr_parameters:delay_nosig_s1_write_n
	wire   [31:0] mm_interconnect_1_nmr_parameters_delay_nosig_s1_writedata;             // mm_interconnect_1:nmr_parameters_delay_nosig_s1_writedata -> nmr_parameters:delay_nosig_s1_writedata
	wire          mm_interconnect_1_nmr_parameters_delay_sig_s1_chipselect;              // mm_interconnect_1:nmr_parameters_delay_sig_s1_chipselect -> nmr_parameters:delay_sig_s1_chipselect
	wire   [31:0] mm_interconnect_1_nmr_parameters_delay_sig_s1_readdata;                // nmr_parameters:delay_sig_s1_readdata -> mm_interconnect_1:nmr_parameters_delay_sig_s1_readdata
	wire    [1:0] mm_interconnect_1_nmr_parameters_delay_sig_s1_address;                 // mm_interconnect_1:nmr_parameters_delay_sig_s1_address -> nmr_parameters:delay_sig_s1_address
	wire          mm_interconnect_1_nmr_parameters_delay_sig_s1_write;                   // mm_interconnect_1:nmr_parameters_delay_sig_s1_write -> nmr_parameters:delay_sig_s1_write_n
	wire   [31:0] mm_interconnect_1_nmr_parameters_delay_sig_s1_writedata;               // mm_interconnect_1:nmr_parameters_delay_sig_s1_writedata -> nmr_parameters:delay_sig_s1_writedata
	wire          mm_interconnect_1_nmr_parameters_delay_t1_s1_chipselect;               // mm_interconnect_1:nmr_parameters_delay_t1_s1_chipselect -> nmr_parameters:delay_t1_s1_chipselect
	wire   [31:0] mm_interconnect_1_nmr_parameters_delay_t1_s1_readdata;                 // nmr_parameters:delay_t1_s1_readdata -> mm_interconnect_1:nmr_parameters_delay_t1_s1_readdata
	wire    [1:0] mm_interconnect_1_nmr_parameters_delay_t1_s1_address;                  // mm_interconnect_1:nmr_parameters_delay_t1_s1_address -> nmr_parameters:delay_t1_s1_address
	wire          mm_interconnect_1_nmr_parameters_delay_t1_s1_write;                    // mm_interconnect_1:nmr_parameters_delay_t1_s1_write -> nmr_parameters:delay_t1_s1_write_n
	wire   [31:0] mm_interconnect_1_nmr_parameters_delay_t1_s1_writedata;                // mm_interconnect_1:nmr_parameters_delay_t1_s1_writedata -> nmr_parameters:delay_t1_s1_writedata
	wire          mm_interconnect_1_nmr_parameters_echoes_per_scan_s1_chipselect;        // mm_interconnect_1:nmr_parameters_echoes_per_scan_s1_chipselect -> nmr_parameters:echoes_per_scan_s1_chipselect
	wire   [31:0] mm_interconnect_1_nmr_parameters_echoes_per_scan_s1_readdata;          // nmr_parameters:echoes_per_scan_s1_readdata -> mm_interconnect_1:nmr_parameters_echoes_per_scan_s1_readdata
	wire    [1:0] mm_interconnect_1_nmr_parameters_echoes_per_scan_s1_address;           // mm_interconnect_1:nmr_parameters_echoes_per_scan_s1_address -> nmr_parameters:echoes_per_scan_s1_address
	wire          mm_interconnect_1_nmr_parameters_echoes_per_scan_s1_write;             // mm_interconnect_1:nmr_parameters_echoes_per_scan_s1_write -> nmr_parameters:echoes_per_scan_s1_write_n
	wire   [31:0] mm_interconnect_1_nmr_parameters_echoes_per_scan_s1_writedata;         // mm_interconnect_1:nmr_parameters_echoes_per_scan_s1_writedata -> nmr_parameters:echoes_per_scan_s1_writedata
	wire   [31:0] mm_interconnect_1_adc_fifo_mem_in_csr_readdata;                        // adc_fifo_mem:wrclk_control_slave_readdata -> mm_interconnect_1:adc_fifo_mem_in_csr_readdata
	wire    [2:0] mm_interconnect_1_adc_fifo_mem_in_csr_address;                         // mm_interconnect_1:adc_fifo_mem_in_csr_address -> adc_fifo_mem:wrclk_control_slave_address
	wire          mm_interconnect_1_adc_fifo_mem_in_csr_read;                            // mm_interconnect_1:adc_fifo_mem_in_csr_read -> adc_fifo_mem:wrclk_control_slave_read
	wire          mm_interconnect_1_adc_fifo_mem_in_csr_write;                           // mm_interconnect_1:adc_fifo_mem_in_csr_write -> adc_fifo_mem:wrclk_control_slave_write
	wire   [31:0] mm_interconnect_1_adc_fifo_mem_in_csr_writedata;                       // mm_interconnect_1:adc_fifo_mem_in_csr_writedata -> adc_fifo_mem:wrclk_control_slave_writedata
	wire   [31:0] mm_interconnect_1_dconv_fifo_mem_in_csr_readdata;                      // dconv_fifo_mem:wrclk_control_slave_readdata -> mm_interconnect_1:dconv_fifo_mem_in_csr_readdata
	wire    [2:0] mm_interconnect_1_dconv_fifo_mem_in_csr_address;                       // mm_interconnect_1:dconv_fifo_mem_in_csr_address -> dconv_fifo_mem:wrclk_control_slave_address
	wire          mm_interconnect_1_dconv_fifo_mem_in_csr_read;                          // mm_interconnect_1:dconv_fifo_mem_in_csr_read -> dconv_fifo_mem:wrclk_control_slave_read
	wire          mm_interconnect_1_dconv_fifo_mem_in_csr_write;                         // mm_interconnect_1:dconv_fifo_mem_in_csr_write -> dconv_fifo_mem:wrclk_control_slave_write
	wire   [31:0] mm_interconnect_1_dconv_fifo_mem_in_csr_writedata;                     // mm_interconnect_1:dconv_fifo_mem_in_csr_writedata -> dconv_fifo_mem:wrclk_control_slave_writedata
	wire   [31:0] mm_interconnect_1_dconv_fifo_mem_q_in_csr_readdata;                    // dconv_fifo_mem_q:wrclk_control_slave_readdata -> mm_interconnect_1:dconv_fifo_mem_q_in_csr_readdata
	wire    [2:0] mm_interconnect_1_dconv_fifo_mem_q_in_csr_address;                     // mm_interconnect_1:dconv_fifo_mem_q_in_csr_address -> dconv_fifo_mem_q:wrclk_control_slave_address
	wire          mm_interconnect_1_dconv_fifo_mem_q_in_csr_read;                        // mm_interconnect_1:dconv_fifo_mem_q_in_csr_read -> dconv_fifo_mem_q:wrclk_control_slave_read
	wire          mm_interconnect_1_dconv_fifo_mem_q_in_csr_write;                       // mm_interconnect_1:dconv_fifo_mem_q_in_csr_write -> dconv_fifo_mem_q:wrclk_control_slave_write
	wire   [31:0] mm_interconnect_1_dconv_fifo_mem_q_in_csr_writedata;                   // mm_interconnect_1:dconv_fifo_mem_q_in_csr_writedata -> dconv_fifo_mem_q:wrclk_control_slave_writedata
	wire          mm_interconnect_1_nmr_parameters_init_delay_s1_chipselect;             // mm_interconnect_1:nmr_parameters_init_delay_s1_chipselect -> nmr_parameters:init_delay_s1_chipselect
	wire   [31:0] mm_interconnect_1_nmr_parameters_init_delay_s1_readdata;               // nmr_parameters:init_delay_s1_readdata -> mm_interconnect_1:nmr_parameters_init_delay_s1_readdata
	wire    [1:0] mm_interconnect_1_nmr_parameters_init_delay_s1_address;                // mm_interconnect_1:nmr_parameters_init_delay_s1_address -> nmr_parameters:init_delay_s1_address
	wire          mm_interconnect_1_nmr_parameters_init_delay_s1_write;                  // mm_interconnect_1:nmr_parameters_init_delay_s1_write -> nmr_parameters:init_delay_s1_write_n
	wire   [31:0] mm_interconnect_1_nmr_parameters_init_delay_s1_writedata;              // mm_interconnect_1:nmr_parameters_init_delay_s1_writedata -> nmr_parameters:init_delay_s1_writedata
	wire   [31:0] mm_interconnect_1_nmr_sys_pll_reconfig_mgmt_avalon_slave_readdata;     // nmr_sys_pll_reconfig:mgmt_readdata -> mm_interconnect_1:nmr_sys_pll_reconfig_mgmt_avalon_slave_readdata
	wire          mm_interconnect_1_nmr_sys_pll_reconfig_mgmt_avalon_slave_waitrequest;  // nmr_sys_pll_reconfig:mgmt_waitrequest -> mm_interconnect_1:nmr_sys_pll_reconfig_mgmt_avalon_slave_waitrequest
	wire    [5:0] mm_interconnect_1_nmr_sys_pll_reconfig_mgmt_avalon_slave_address;      // mm_interconnect_1:nmr_sys_pll_reconfig_mgmt_avalon_slave_address -> nmr_sys_pll_reconfig:mgmt_address
	wire          mm_interconnect_1_nmr_sys_pll_reconfig_mgmt_avalon_slave_read;         // mm_interconnect_1:nmr_sys_pll_reconfig_mgmt_avalon_slave_read -> nmr_sys_pll_reconfig:mgmt_read
	wire          mm_interconnect_1_nmr_sys_pll_reconfig_mgmt_avalon_slave_write;        // mm_interconnect_1:nmr_sys_pll_reconfig_mgmt_avalon_slave_write -> nmr_sys_pll_reconfig:mgmt_write
	wire   [31:0] mm_interconnect_1_nmr_sys_pll_reconfig_mgmt_avalon_slave_writedata;    // mm_interconnect_1:nmr_sys_pll_reconfig_mgmt_avalon_slave_writedata -> nmr_sys_pll_reconfig:mgmt_writedata
	wire   [31:0] mm_interconnect_1_analyzer_pll_reconfig_mgmt_avalon_slave_readdata;    // analyzer_pll_reconfig:mgmt_readdata -> mm_interconnect_1:analyzer_pll_reconfig_mgmt_avalon_slave_readdata
	wire          mm_interconnect_1_analyzer_pll_reconfig_mgmt_avalon_slave_waitrequest; // analyzer_pll_reconfig:mgmt_waitrequest -> mm_interconnect_1:analyzer_pll_reconfig_mgmt_avalon_slave_waitrequest
	wire    [5:0] mm_interconnect_1_analyzer_pll_reconfig_mgmt_avalon_slave_address;     // mm_interconnect_1:analyzer_pll_reconfig_mgmt_avalon_slave_address -> analyzer_pll_reconfig:mgmt_address
	wire          mm_interconnect_1_analyzer_pll_reconfig_mgmt_avalon_slave_read;        // mm_interconnect_1:analyzer_pll_reconfig_mgmt_avalon_slave_read -> analyzer_pll_reconfig:mgmt_read
	wire          mm_interconnect_1_analyzer_pll_reconfig_mgmt_avalon_slave_write;       // mm_interconnect_1:analyzer_pll_reconfig_mgmt_avalon_slave_write -> analyzer_pll_reconfig:mgmt_write
	wire   [31:0] mm_interconnect_1_analyzer_pll_reconfig_mgmt_avalon_slave_writedata;   // mm_interconnect_1:analyzer_pll_reconfig_mgmt_avalon_slave_writedata -> analyzer_pll_reconfig:mgmt_writedata
	wire   [31:0] mm_interconnect_1_dconv_fifo_mem_out_readdata;                         // dconv_fifo_mem:avalonmm_read_slave_readdata -> mm_interconnect_1:dconv_fifo_mem_out_readdata
	wire          mm_interconnect_1_dconv_fifo_mem_out_waitrequest;                      // dconv_fifo_mem:avalonmm_read_slave_waitrequest -> mm_interconnect_1:dconv_fifo_mem_out_waitrequest
	wire    [0:0] mm_interconnect_1_dconv_fifo_mem_out_address;                          // mm_interconnect_1:dconv_fifo_mem_out_address -> dconv_fifo_mem:avalonmm_read_slave_address
	wire          mm_interconnect_1_dconv_fifo_mem_out_read;                             // mm_interconnect_1:dconv_fifo_mem_out_read -> dconv_fifo_mem:avalonmm_read_slave_read
	wire   [31:0] mm_interconnect_1_dconv_fifo_mem_q_out_readdata;                       // dconv_fifo_mem_q:avalonmm_read_slave_readdata -> mm_interconnect_1:dconv_fifo_mem_q_out_readdata
	wire          mm_interconnect_1_dconv_fifo_mem_q_out_waitrequest;                    // dconv_fifo_mem_q:avalonmm_read_slave_waitrequest -> mm_interconnect_1:dconv_fifo_mem_q_out_waitrequest
	wire    [0:0] mm_interconnect_1_dconv_fifo_mem_q_out_address;                        // mm_interconnect_1:dconv_fifo_mem_q_out_address -> dconv_fifo_mem_q:avalonmm_read_slave_address
	wire          mm_interconnect_1_dconv_fifo_mem_q_out_read;                           // mm_interconnect_1:dconv_fifo_mem_q_out_read -> dconv_fifo_mem_q:avalonmm_read_slave_read
	wire          mm_interconnect_1_nmr_parameters_pulse_180deg_s1_chipselect;           // mm_interconnect_1:nmr_parameters_pulse_180deg_s1_chipselect -> nmr_parameters:pulse_180deg_s1_chipselect
	wire   [31:0] mm_interconnect_1_nmr_parameters_pulse_180deg_s1_readdata;             // nmr_parameters:pulse_180deg_s1_readdata -> mm_interconnect_1:nmr_parameters_pulse_180deg_s1_readdata
	wire    [1:0] mm_interconnect_1_nmr_parameters_pulse_180deg_s1_address;              // mm_interconnect_1:nmr_parameters_pulse_180deg_s1_address -> nmr_parameters:pulse_180deg_s1_address
	wire          mm_interconnect_1_nmr_parameters_pulse_180deg_s1_write;                // mm_interconnect_1:nmr_parameters_pulse_180deg_s1_write -> nmr_parameters:pulse_180deg_s1_write_n
	wire   [31:0] mm_interconnect_1_nmr_parameters_pulse_180deg_s1_writedata;            // mm_interconnect_1:nmr_parameters_pulse_180deg_s1_writedata -> nmr_parameters:pulse_180deg_s1_writedata
	wire          mm_interconnect_1_nmr_parameters_pulse_90deg_s1_chipselect;            // mm_interconnect_1:nmr_parameters_pulse_90deg_s1_chipselect -> nmr_parameters:pulse_90deg_s1_chipselect
	wire   [31:0] mm_interconnect_1_nmr_parameters_pulse_90deg_s1_readdata;              // nmr_parameters:pulse_90deg_s1_readdata -> mm_interconnect_1:nmr_parameters_pulse_90deg_s1_readdata
	wire    [1:0] mm_interconnect_1_nmr_parameters_pulse_90deg_s1_address;               // mm_interconnect_1:nmr_parameters_pulse_90deg_s1_address -> nmr_parameters:pulse_90deg_s1_address
	wire          mm_interconnect_1_nmr_parameters_pulse_90deg_s1_write;                 // mm_interconnect_1:nmr_parameters_pulse_90deg_s1_write -> nmr_parameters:pulse_90deg_s1_write_n
	wire   [31:0] mm_interconnect_1_nmr_parameters_pulse_90deg_s1_writedata;             // mm_interconnect_1:nmr_parameters_pulse_90deg_s1_writedata -> nmr_parameters:pulse_90deg_s1_writedata
	wire          mm_interconnect_1_nmr_parameters_pulse_t1_s1_chipselect;               // mm_interconnect_1:nmr_parameters_pulse_t1_s1_chipselect -> nmr_parameters:pulse_t1_s1_chipselect
	wire   [31:0] mm_interconnect_1_nmr_parameters_pulse_t1_s1_readdata;                 // nmr_parameters:pulse_t1_s1_readdata -> mm_interconnect_1:nmr_parameters_pulse_t1_s1_readdata
	wire    [1:0] mm_interconnect_1_nmr_parameters_pulse_t1_s1_address;                  // mm_interconnect_1:nmr_parameters_pulse_t1_s1_address -> nmr_parameters:pulse_t1_s1_address
	wire          mm_interconnect_1_nmr_parameters_pulse_t1_s1_write;                    // mm_interconnect_1:nmr_parameters_pulse_t1_s1_write -> nmr_parameters:pulse_t1_s1_write_n
	wire   [31:0] mm_interconnect_1_nmr_parameters_pulse_t1_s1_writedata;                // mm_interconnect_1:nmr_parameters_pulse_t1_s1_writedata -> nmr_parameters:pulse_t1_s1_writedata
	wire          mm_interconnect_1_nmr_parameters_rx_delay_s1_chipselect;               // mm_interconnect_1:nmr_parameters_rx_delay_s1_chipselect -> nmr_parameters:rx_delay_s1_chipselect
	wire   [31:0] mm_interconnect_1_nmr_parameters_rx_delay_s1_readdata;                 // nmr_parameters:rx_delay_s1_readdata -> mm_interconnect_1:nmr_parameters_rx_delay_s1_readdata
	wire    [1:0] mm_interconnect_1_nmr_parameters_rx_delay_s1_address;                  // mm_interconnect_1:nmr_parameters_rx_delay_s1_address -> nmr_parameters:rx_delay_s1_address
	wire          mm_interconnect_1_nmr_parameters_rx_delay_s1_write;                    // mm_interconnect_1:nmr_parameters_rx_delay_s1_write -> nmr_parameters:rx_delay_s1_write_n
	wire   [31:0] mm_interconnect_1_nmr_parameters_rx_delay_s1_writedata;                // mm_interconnect_1:nmr_parameters_rx_delay_s1_writedata -> nmr_parameters:rx_delay_s1_writedata
	wire          mm_interconnect_1_ctrl_out_s1_chipselect;                              // mm_interconnect_1:ctrl_out_s1_chipselect -> ctrl_out:chipselect
	wire   [31:0] mm_interconnect_1_ctrl_out_s1_readdata;                                // ctrl_out:readdata -> mm_interconnect_1:ctrl_out_s1_readdata
	wire    [1:0] mm_interconnect_1_ctrl_out_s1_address;                                 // mm_interconnect_1:ctrl_out_s1_address -> ctrl_out:address
	wire          mm_interconnect_1_ctrl_out_s1_write;                                   // mm_interconnect_1:ctrl_out_s1_write -> ctrl_out:write_n
	wire   [31:0] mm_interconnect_1_ctrl_out_s1_writedata;                               // mm_interconnect_1:ctrl_out_s1_writedata -> ctrl_out:writedata
	wire   [31:0] mm_interconnect_1_ctrl_in_s1_readdata;                                 // ctrl_in:readdata -> mm_interconnect_1:ctrl_in_s1_readdata
	wire    [1:0] mm_interconnect_1_ctrl_in_s1_address;                                  // mm_interconnect_1:ctrl_in_s1_address -> ctrl_in:address
	wire          mm_interconnect_1_aux_cnt_out_s1_chipselect;                           // mm_interconnect_1:aux_cnt_out_s1_chipselect -> aux_cnt_out:chipselect
	wire   [31:0] mm_interconnect_1_aux_cnt_out_s1_readdata;                             // aux_cnt_out:readdata -> mm_interconnect_1:aux_cnt_out_s1_readdata
	wire    [1:0] mm_interconnect_1_aux_cnt_out_s1_address;                              // mm_interconnect_1:aux_cnt_out_s1_address -> aux_cnt_out:address
	wire          mm_interconnect_1_aux_cnt_out_s1_write;                                // mm_interconnect_1:aux_cnt_out_s1_write -> aux_cnt_out:write_n
	wire   [31:0] mm_interconnect_1_aux_cnt_out_s1_writedata;                            // mm_interconnect_1:aux_cnt_out_s1_writedata -> aux_cnt_out:writedata
	wire          mm_interconnect_1_nmr_parameters_samples_per_echo_s1_chipselect;       // mm_interconnect_1:nmr_parameters_samples_per_echo_s1_chipselect -> nmr_parameters:samples_per_echo_s1_chipselect
	wire   [31:0] mm_interconnect_1_nmr_parameters_samples_per_echo_s1_readdata;         // nmr_parameters:samples_per_echo_s1_readdata -> mm_interconnect_1:nmr_parameters_samples_per_echo_s1_readdata
	wire    [1:0] mm_interconnect_1_nmr_parameters_samples_per_echo_s1_address;          // mm_interconnect_1:nmr_parameters_samples_per_echo_s1_address -> nmr_parameters:samples_per_echo_s1_address
	wire          mm_interconnect_1_nmr_parameters_samples_per_echo_s1_write;            // mm_interconnect_1:nmr_parameters_samples_per_echo_s1_write -> nmr_parameters:samples_per_echo_s1_write_n
	wire   [31:0] mm_interconnect_1_nmr_parameters_samples_per_echo_s1_writedata;        // mm_interconnect_1:nmr_parameters_samples_per_echo_s1_writedata -> nmr_parameters:samples_per_echo_s1_writedata
	wire          mm_interconnect_1_dac_grad_spi_control_port_chipselect;                // mm_interconnect_1:dac_grad_spi_control_port_chipselect -> dac_grad:spi_select
	wire   [31:0] mm_interconnect_1_dac_grad_spi_control_port_readdata;                  // dac_grad:data_to_cpu -> mm_interconnect_1:dac_grad_spi_control_port_readdata
	wire    [2:0] mm_interconnect_1_dac_grad_spi_control_port_address;                   // mm_interconnect_1:dac_grad_spi_control_port_address -> dac_grad:mem_addr
	wire          mm_interconnect_1_dac_grad_spi_control_port_read;                      // mm_interconnect_1:dac_grad_spi_control_port_read -> dac_grad:read_n
	wire          mm_interconnect_1_dac_grad_spi_control_port_write;                     // mm_interconnect_1:dac_grad_spi_control_port_write -> dac_grad:write_n
	wire   [31:0] mm_interconnect_1_dac_grad_spi_control_port_writedata;                 // mm_interconnect_1:dac_grad_spi_control_port_writedata -> dac_grad:data_from_cpu
	wire          mm_interconnect_1_spi_mtch_ntwrk_spi_control_port_chipselect;          // mm_interconnect_1:spi_mtch_ntwrk_spi_control_port_chipselect -> spi_mtch_ntwrk:spi_select
	wire   [31:0] mm_interconnect_1_spi_mtch_ntwrk_spi_control_port_readdata;            // spi_mtch_ntwrk:data_to_cpu -> mm_interconnect_1:spi_mtch_ntwrk_spi_control_port_readdata
	wire    [2:0] mm_interconnect_1_spi_mtch_ntwrk_spi_control_port_address;             // mm_interconnect_1:spi_mtch_ntwrk_spi_control_port_address -> spi_mtch_ntwrk:mem_addr
	wire          mm_interconnect_1_spi_mtch_ntwrk_spi_control_port_read;                // mm_interconnect_1:spi_mtch_ntwrk_spi_control_port_read -> spi_mtch_ntwrk:read_n
	wire          mm_interconnect_1_spi_mtch_ntwrk_spi_control_port_write;               // mm_interconnect_1:spi_mtch_ntwrk_spi_control_port_write -> spi_mtch_ntwrk:write_n
	wire   [31:0] mm_interconnect_1_spi_mtch_ntwrk_spi_control_port_writedata;           // mm_interconnect_1:spi_mtch_ntwrk_spi_control_port_writedata -> spi_mtch_ntwrk:data_from_cpu
	wire          mm_interconnect_1_spi_afe_relays_spi_control_port_chipselect;          // mm_interconnect_1:spi_afe_relays_spi_control_port_chipselect -> spi_afe_relays:spi_select
	wire   [31:0] mm_interconnect_1_spi_afe_relays_spi_control_port_readdata;            // spi_afe_relays:data_to_cpu -> mm_interconnect_1:spi_afe_relays_spi_control_port_readdata
	wire    [2:0] mm_interconnect_1_spi_afe_relays_spi_control_port_address;             // mm_interconnect_1:spi_afe_relays_spi_control_port_address -> spi_afe_relays:mem_addr
	wire          mm_interconnect_1_spi_afe_relays_spi_control_port_read;                // mm_interconnect_1:spi_afe_relays_spi_control_port_read -> spi_afe_relays:read_n
	wire          mm_interconnect_1_spi_afe_relays_spi_control_port_write;               // mm_interconnect_1:spi_afe_relays_spi_control_port_write -> spi_afe_relays:write_n
	wire   [31:0] mm_interconnect_1_spi_afe_relays_spi_control_port_writedata;           // mm_interconnect_1:spi_afe_relays_spi_control_port_writedata -> spi_afe_relays:data_from_cpu
	wire          mm_interconnect_1_dma_fifo_control_port_slave_chipselect;              // mm_interconnect_1:dma_fifo_control_port_slave_chipselect -> dma_fifo:dma_ctl_chipselect
	wire   [31:0] mm_interconnect_1_dma_fifo_control_port_slave_readdata;                // dma_fifo:dma_ctl_readdata -> mm_interconnect_1:dma_fifo_control_port_slave_readdata
	wire    [2:0] mm_interconnect_1_dma_fifo_control_port_slave_address;                 // mm_interconnect_1:dma_fifo_control_port_slave_address -> dma_fifo:dma_ctl_address
	wire          mm_interconnect_1_dma_fifo_control_port_slave_write;                   // mm_interconnect_1:dma_fifo_control_port_slave_write -> dma_fifo:dma_ctl_write_n
	wire   [31:0] mm_interconnect_1_dma_fifo_control_port_slave_writedata;               // mm_interconnect_1:dma_fifo_control_port_slave_writedata -> dma_fifo:dma_ctl_writedata
	wire          mm_interconnect_1_dma_dconvi_control_port_slave_chipselect;            // mm_interconnect_1:dma_dconvi_control_port_slave_chipselect -> dma_dconvi:dma_ctl_chipselect
	wire   [31:0] mm_interconnect_1_dma_dconvi_control_port_slave_readdata;              // dma_dconvi:dma_ctl_readdata -> mm_interconnect_1:dma_dconvi_control_port_slave_readdata
	wire    [2:0] mm_interconnect_1_dma_dconvi_control_port_slave_address;               // mm_interconnect_1:dma_dconvi_control_port_slave_address -> dma_dconvi:dma_ctl_address
	wire          mm_interconnect_1_dma_dconvi_control_port_slave_write;                 // mm_interconnect_1:dma_dconvi_control_port_slave_write -> dma_dconvi:dma_ctl_write_n
	wire   [31:0] mm_interconnect_1_dma_dconvi_control_port_slave_writedata;             // mm_interconnect_1:dma_dconvi_control_port_slave_writedata -> dma_dconvi:dma_ctl_writedata
	wire          mm_interconnect_1_dma_dconvq_control_port_slave_chipselect;            // mm_interconnect_1:dma_dconvq_control_port_slave_chipselect -> dma_dconvq:dma_ctl_chipselect
	wire   [31:0] mm_interconnect_1_dma_dconvq_control_port_slave_readdata;              // dma_dconvq:dma_ctl_readdata -> mm_interconnect_1:dma_dconvq_control_port_slave_readdata
	wire    [2:0] mm_interconnect_1_dma_dconvq_control_port_slave_address;               // mm_interconnect_1:dma_dconvq_control_port_slave_address -> dma_dconvq:dma_ctl_address
	wire          mm_interconnect_1_dma_dconvq_control_port_slave_write;                 // mm_interconnect_1:dma_dconvq_control_port_slave_write -> dma_dconvq:dma_ctl_write_n
	wire   [31:0] mm_interconnect_1_dma_dconvq_control_port_slave_writedata;             // mm_interconnect_1:dma_dconvq_control_port_slave_writedata -> dma_dconvq:dma_ctl_writedata
	wire          mm_interconnect_1_dma_dummy_control_port_slave_chipselect;             // mm_interconnect_1:dma_dummy_control_port_slave_chipselect -> dma_dummy:dma_ctl_chipselect
	wire   [31:0] mm_interconnect_1_dma_dummy_control_port_slave_readdata;               // dma_dummy:dma_ctl_readdata -> mm_interconnect_1:dma_dummy_control_port_slave_readdata
	wire    [2:0] mm_interconnect_1_dma_dummy_control_port_slave_address;                // mm_interconnect_1:dma_dummy_control_port_slave_address -> dma_dummy:dma_ctl_address
	wire          mm_interconnect_1_dma_dummy_control_port_slave_write;                  // mm_interconnect_1:dma_dummy_control_port_slave_write -> dma_dummy:dma_ctl_write_n
	wire   [31:0] mm_interconnect_1_dma_dummy_control_port_slave_writedata;              // mm_interconnect_1:dma_dummy_control_port_slave_writedata -> dma_dummy:dma_ctl_writedata
	wire          irq_mapper_receiver0_irq;                                              // alt_vip_vfr_vga:slave_irq -> irq_mapper:receiver0_irq
	wire          irq_mapper_receiver1_irq;                                              // jtag_uart:av_irq -> irq_mapper:receiver1_irq
	wire   [31:0] hps_0_f2h_irq0_irq;                                                    // irq_mapper:sender_irq -> hps_0:f2h_irq_p0
	wire          irq_mapper_001_receiver0_irq;                                          // i2c_int:intr -> irq_mapper_001:receiver0_irq
	wire          irq_mapper_001_receiver1_irq;                                          // i2c_ext:intr -> irq_mapper_001:receiver1_irq
	wire          irq_mapper_001_receiver2_irq;                                          // dac_grad:irq -> irq_mapper_001:receiver2_irq
	wire          irq_mapper_001_receiver3_irq;                                          // dma_fifo:dma_ctl_irq -> irq_mapper_001:receiver3_irq
	wire          irq_mapper_001_receiver4_irq;                                          // spi_mtch_ntwrk:irq -> irq_mapper_001:receiver4_irq
	wire          irq_mapper_001_receiver5_irq;                                          // dma_dconvi:dma_ctl_irq -> irq_mapper_001:receiver5_irq
	wire          irq_mapper_001_receiver6_irq;                                          // dma_dconvq:dma_ctl_irq -> irq_mapper_001:receiver6_irq
	wire          irq_mapper_001_receiver7_irq;                                          // spi_afe_relays:irq -> irq_mapper_001:receiver7_irq
	wire   [31:0] hps_0_f2h_irq1_irq;                                                    // irq_mapper_001:sender_irq -> hps_0:f2h_irq_p1
	wire          adc_fifo_dc_out_valid;                                                 // adc_fifo_dc:out_valid -> avalon_st_adapter:in_0_valid
	wire   [15:0] adc_fifo_dc_out_data;                                                  // adc_fifo_dc:out_data -> avalon_st_adapter:in_0_data
	wire          adc_fifo_dc_out_ready;                                                 // avalon_st_adapter:in_0_ready -> adc_fifo_dc:out_ready
	wire          avalon_st_adapter_out_0_valid;                                         // avalon_st_adapter:out_0_valid -> adc_fifo_mem:avalonst_sink_valid
	wire   [31:0] avalon_st_adapter_out_0_data;                                          // avalon_st_adapter:out_0_data -> adc_fifo_mem:avalonst_sink_data
	wire          avalon_st_adapter_out_0_ready;                                         // adc_fifo_mem:avalonst_sink_ready -> avalon_st_adapter:out_0_ready
	wire          dconv_fifo_dc_out_valid;                                               // dconv_fifo_dc:out_valid -> avalon_st_adapter_001:in_0_valid
	wire   [31:0] dconv_fifo_dc_out_data;                                                // dconv_fifo_dc:out_data -> avalon_st_adapter_001:in_0_data
	wire          dconv_fifo_dc_out_ready;                                               // avalon_st_adapter_001:in_0_ready -> dconv_fifo_dc:out_ready
	wire          avalon_st_adapter_001_out_0_valid;                                     // avalon_st_adapter_001:out_0_valid -> dconv_fifo_mem:avalonst_sink_valid
	wire   [31:0] avalon_st_adapter_001_out_0_data;                                      // avalon_st_adapter_001:out_0_data -> dconv_fifo_mem:avalonst_sink_data
	wire          avalon_st_adapter_001_out_0_ready;                                     // dconv_fifo_mem:avalonst_sink_ready -> avalon_st_adapter_001:out_0_ready
	wire          dconv_fifo_dc_q_out_valid;                                             // dconv_fifo_dc_q:out_valid -> avalon_st_adapter_002:in_0_valid
	wire   [31:0] dconv_fifo_dc_q_out_data;                                              // dconv_fifo_dc_q:out_data -> avalon_st_adapter_002:in_0_data
	wire          dconv_fifo_dc_q_out_ready;                                             // avalon_st_adapter_002:in_0_ready -> dconv_fifo_dc_q:out_ready
	wire          avalon_st_adapter_002_out_0_valid;                                     // avalon_st_adapter_002:out_0_valid -> dconv_fifo_mem_q:avalonst_sink_valid
	wire   [31:0] avalon_st_adapter_002_out_0_data;                                      // avalon_st_adapter_002:out_0_data -> dconv_fifo_mem_q:avalonst_sink_data
	wire          avalon_st_adapter_002_out_0_ready;                                     // dconv_fifo_mem_q:avalonst_sink_ready -> avalon_st_adapter_002:out_0_ready
	wire          rst_controller_reset_out_reset;                                        // rst_controller:reset_out -> [adc_fifo_dc:in_reset_n, dconv_fifo_dc:in_reset_n, dconv_fifo_dc_q:in_reset_n]
	wire          rst_controller_001_reset_out_reset;                                    // rst_controller_001:reset_out -> [adc_fifo_dc:out_reset_n, adc_fifo_mem:reset_n, avalon_st_adapter:in_rst_0_reset, avalon_st_adapter_001:in_rst_0_reset, avalon_st_adapter_002:in_rst_0_reset, dconv_fifo_dc:out_reset_n, dconv_fifo_dc_q:out_reset_n, dconv_fifo_mem:reset_n, dconv_fifo_mem_q:reset_n, mm_interconnect_1:adc_fifo_mem_reset_in_reset_bridge_in_reset_reset]
	wire          rst_controller_002_reset_out_reset;                                    // rst_controller_002:reset_out -> [alt_vip_itc_0:rst, alt_vip_vfr_vga:reset, mm_interconnect_1:alt_vip_vfr_vga_clock_reset_reset_reset_bridge_in_reset_reset]
	wire          rst_controller_003_reset_out_reset;                                    // rst_controller_003:reset_out -> [alt_vip_vfr_vga:master_reset, analyzer_pll_reconfig:mgmt_reset, aux_cnt_out:reset_n, ctrl_in:reset_n, ctrl_out:reset_n, dac_grad:reset_n, dconv_fir:coeff_in_areset, dconv_fir_q:coeff_in_areset, dma_dconvi:system_reset_n, dma_dconvq:system_reset_n, dma_dummy:system_reset_n, dma_fifo:system_reset_n, fifo_dummy64_in:reset_n, fifo_dummy64_out:reset_n, fifo_dummy:reset_n, i2c_ext:rst_n, i2c_int:rst_n, jtag_uart:rst_n, mm_interconnect_0:alt_vip_vfr_vga_clock_master_reset_reset_bridge_in_reset_reset, mm_interconnect_0:master_secure_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_1:dma_fifo_reset_reset_bridge_in_reset_reset, mm_interconnect_1:master_non_sec_clk_reset_reset_bridge_in_reset_reset, nmr_parameters:adc_val_sub_reset_reset_n, nmr_parameters:delay_nosig_reset_reset_n, nmr_parameters:delay_sig_reset_reset_n, nmr_parameters:delay_t1_reset_reset_n, nmr_parameters:echoes_per_scan_reset_reset_n, nmr_parameters:init_delay_reset_reset_n, nmr_parameters:pulse_180deg_reset_reset_n, nmr_parameters:pulse_90deg_reset_reset_n, nmr_parameters:pulse_t1_reset_reset_n, nmr_parameters:rx_delay_reset_reset_n, nmr_parameters:samples_per_echo_reset_reset_n, nmr_sys_pll_reconfig:mgmt_reset, sdram:reset_n, spi_afe_relays:reset_n, spi_mtch_ntwrk:reset_n, switches:reset_n, sysid_qsys:reset_n]
	wire          rst_controller_004_reset_out_reset;                                    // rst_controller_004:reset_out -> [mm_interconnect_0:hps_0_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_1:hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset]

	altera_avalon_dc_fifo #(
		.SYMBOLS_PER_BEAT   (1),
		.BITS_PER_SYMBOL    (16),
		.FIFO_DEPTH         (16384),
		.CHANNEL_WIDTH      (0),
		.ERROR_WIDTH        (0),
		.USE_PACKETS        (0),
		.USE_IN_FILL_LEVEL  (0),
		.USE_OUT_FILL_LEVEL (0),
		.WR_SYNC_DEPTH      (3),
		.RD_SYNC_DEPTH      (3)
	) adc_fifo_dc (
		.in_clk            (fifo_clk_bridge_in_clk),               //        in_clk.clk
		.in_reset_n        (~rst_controller_reset_out_reset),      //  in_clk_reset.reset_n
		.out_clk           (clk_clk),                              //       out_clk.clk
		.out_reset_n       (~rst_controller_001_reset_out_reset),  // out_clk_reset.reset_n
		.in_data           (adc_fifo_in_data),                     //            in.data
		.in_valid          (adc_fifo_in_valid),                    //              .valid
		.in_ready          (adc_fifo_in_ready),                    //              .ready
		.out_data          (adc_fifo_dc_out_data),                 //           out.data
		.out_valid         (adc_fifo_dc_out_valid),                //              .valid
		.out_ready         (adc_fifo_dc_out_ready),                //              .ready
		.in_csr_address    (1'b0),                                 //   (terminated)
		.in_csr_read       (1'b0),                                 //   (terminated)
		.in_csr_write      (1'b0),                                 //   (terminated)
		.in_csr_readdata   (),                                     //   (terminated)
		.in_csr_writedata  (32'b00000000000000000000000000000000), //   (terminated)
		.out_csr_address   (1'b0),                                 //   (terminated)
		.out_csr_read      (1'b0),                                 //   (terminated)
		.out_csr_write     (1'b0),                                 //   (terminated)
		.out_csr_readdata  (),                                     //   (terminated)
		.out_csr_writedata (32'b00000000000000000000000000000000), //   (terminated)
		.in_startofpacket  (1'b0),                                 //   (terminated)
		.in_endofpacket    (1'b0),                                 //   (terminated)
		.out_startofpacket (),                                     //   (terminated)
		.out_endofpacket   (),                                     //   (terminated)
		.in_empty          (1'b0),                                 //   (terminated)
		.out_empty         (),                                     //   (terminated)
		.in_error          (1'b0),                                 //   (terminated)
		.out_error         (),                                     //   (terminated)
		.in_channel        (1'b0),                                 //   (terminated)
		.out_channel       (),                                     //   (terminated)
		.space_avail_data  ()                                      //   (terminated)
	);

	soc_system_v5_adc_fifo_mem adc_fifo_mem (
		.wrclock                         (clk_clk),                                         //   clk_in.clk
		.reset_n                         (~rst_controller_001_reset_out_reset),             // reset_in.reset_n
		.avalonst_sink_valid             (avalon_st_adapter_out_0_valid),                   //       in.valid
		.avalonst_sink_data              (avalon_st_adapter_out_0_data),                    //         .data
		.avalonst_sink_ready             (avalon_st_adapter_out_0_ready),                   //         .ready
		.avalonmm_read_slave_readdata    (mm_interconnect_1_adc_fifo_mem_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read        (mm_interconnect_1_adc_fifo_mem_out_read),         //         .read
		.avalonmm_read_slave_address     (mm_interconnect_1_adc_fifo_mem_out_address),      //         .address
		.avalonmm_read_slave_waitrequest (mm_interconnect_1_adc_fifo_mem_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address     (mm_interconnect_1_adc_fifo_mem_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read        (mm_interconnect_1_adc_fifo_mem_in_csr_read),      //         .read
		.wrclk_control_slave_writedata   (mm_interconnect_1_adc_fifo_mem_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write       (mm_interconnect_1_adc_fifo_mem_in_csr_write),     //         .write
		.wrclk_control_slave_readdata    (mm_interconnect_1_adc_fifo_mem_in_csr_readdata)   //         .readdata
	);

	alt_vipitc131_IS2Vid #(
		.NUMBER_OF_COLOUR_PLANES       (4),
		.COLOUR_PLANES_ARE_IN_PARALLEL (1),
		.BPS                           (8),
		.INTERLACED                    (0),
		.H_ACTIVE_PIXELS               (1024),
		.V_ACTIVE_LINES                (768),
		.ACCEPT_COLOURS_IN_SEQ         (0),
		.FIFO_DEPTH                    (1920),
		.CLOCKS_ARE_SAME               (0),
		.USE_CONTROL                   (0),
		.NO_OF_MODES                   (1),
		.THRESHOLD                     (1919),
		.STD_WIDTH                     (1),
		.GENERATE_SYNC                 (0),
		.USE_EMBEDDED_SYNCS            (0),
		.AP_LINE                       (0),
		.V_BLANK                       (0),
		.H_BLANK                       (0),
		.H_SYNC_LENGTH                 (136),
		.H_FRONT_PORCH                 (24),
		.H_BACK_PORCH                  (160),
		.V_SYNC_LENGTH                 (6),
		.V_FRONT_PORCH                 (3),
		.V_BACK_PORCH                  (29),
		.F_RISING_EDGE                 (0),
		.F_FALLING_EDGE                (0),
		.FIELD0_V_RISING_EDGE          (0),
		.FIELD0_V_BLANK                (0),
		.FIELD0_V_SYNC_LENGTH          (0),
		.FIELD0_V_FRONT_PORCH          (0),
		.FIELD0_V_BACK_PORCH           (0),
		.ANC_LINE                      (0),
		.FIELD0_ANC_LINE               (0)
	) alt_vip_itc_0 (
		.is_clk        (gp_pll_outclk0_clk),                                    //       is_clk_rst.clk
		.rst           (rst_controller_002_reset_out_reset),                    // is_clk_rst_reset.reset
		.is_data       (alt_vip_vfr_vga_avalon_streaming_source_data),          //              din.data
		.is_valid      (alt_vip_vfr_vga_avalon_streaming_source_valid),         //                 .valid
		.is_ready      (alt_vip_vfr_vga_avalon_streaming_source_ready),         //                 .ready
		.is_sop        (alt_vip_vfr_vga_avalon_streaming_source_startofpacket), //                 .startofpacket
		.is_eop        (alt_vip_vfr_vga_avalon_streaming_source_endofpacket),   //                 .endofpacket
		.vid_clk       (alt_vip_itc_0_clocked_video_vid_clk),                   //    clocked_video.export
		.vid_data      (alt_vip_itc_0_clocked_video_vid_data),                  //                 .export
		.underflow     (alt_vip_itc_0_clocked_video_underflow),                 //                 .export
		.vid_datavalid (alt_vip_itc_0_clocked_video_vid_datavalid),             //                 .export
		.vid_v_sync    (alt_vip_itc_0_clocked_video_vid_v_sync),                //                 .export
		.vid_h_sync    (alt_vip_itc_0_clocked_video_vid_h_sync),                //                 .export
		.vid_f         (alt_vip_itc_0_clocked_video_vid_f),                     //                 .export
		.vid_h         (alt_vip_itc_0_clocked_video_vid_h),                     //                 .export
		.vid_v         (alt_vip_itc_0_clocked_video_vid_v)                      //                 .export
	);

	alt_vipvfr131_vfr #(
		.BITS_PER_PIXEL_PER_COLOR_PLANE (8),
		.NUMBER_OF_CHANNELS_IN_PARALLEL (4),
		.NUMBER_OF_CHANNELS_IN_SEQUENCE (1),
		.MAX_IMAGE_WIDTH                (1024),
		.MAX_IMAGE_HEIGHT               (768),
		.MEM_PORT_WIDTH                 (128),
		.RMASTER_FIFO_DEPTH             (64),
		.RMASTER_BURST_TARGET           (32),
		.CLOCKS_ARE_SEPARATE            (1)
	) alt_vip_vfr_vga (
		.clock                (gp_pll_outclk0_clk),                                       //             clock_reset.clk
		.reset                (rst_controller_002_reset_out_reset),                       //       clock_reset_reset.reset
		.master_clock         (clk_clk),                                                  //            clock_master.clk
		.master_reset         (rst_controller_003_reset_out_reset),                       //      clock_master_reset.reset
		.slave_address        (mm_interconnect_1_alt_vip_vfr_vga_avalon_slave_address),   //            avalon_slave.address
		.slave_write          (mm_interconnect_1_alt_vip_vfr_vga_avalon_slave_write),     //                        .write
		.slave_writedata      (mm_interconnect_1_alt_vip_vfr_vga_avalon_slave_writedata), //                        .writedata
		.slave_read           (mm_interconnect_1_alt_vip_vfr_vga_avalon_slave_read),      //                        .read
		.slave_readdata       (mm_interconnect_1_alt_vip_vfr_vga_avalon_slave_readdata),  //                        .readdata
		.slave_irq            (irq_mapper_receiver0_irq),                                 //        interrupt_sender.irq
		.dout_data            (alt_vip_vfr_vga_avalon_streaming_source_data),             // avalon_streaming_source.data
		.dout_valid           (alt_vip_vfr_vga_avalon_streaming_source_valid),            //                        .valid
		.dout_ready           (alt_vip_vfr_vga_avalon_streaming_source_ready),            //                        .ready
		.dout_startofpacket   (alt_vip_vfr_vga_avalon_streaming_source_startofpacket),    //                        .startofpacket
		.dout_endofpacket     (alt_vip_vfr_vga_avalon_streaming_source_endofpacket),      //                        .endofpacket
		.master_address       (alt_vip_vfr_vga_avalon_master_address),                    //           avalon_master.address
		.master_burstcount    (alt_vip_vfr_vga_avalon_master_burstcount),                 //                        .burstcount
		.master_readdata      (alt_vip_vfr_vga_avalon_master_readdata),                   //                        .readdata
		.master_read          (alt_vip_vfr_vga_avalon_master_read),                       //                        .read
		.master_readdatavalid (alt_vip_vfr_vga_avalon_master_readdatavalid),              //                        .readdatavalid
		.master_waitrequest   (alt_vip_vfr_vga_avalon_master_waitrequest)                 //                        .waitrequest
	);

	soc_system_v5_analyzer_pll analyzer_pll (
		.refclk            (clk_clk),                                               //            refclk.clk
		.rst               (analyzer_pll_reset_reset),                              //             reset.reset
		.outclk_0          (analyzer_pll_outclk0_clk),                              //           outclk0.clk
		.outclk_1          (analyzer_pll_outclk1_clk),                              //           outclk1.clk
		.outclk_2          (analyzer_pll_outclk2_clk),                              //           outclk2.clk
		.outclk_3          (analyzer_pll_outclk3_clk),                              //           outclk3.clk
		.locked            (analyzer_pll_locked_export),                            //            locked.export
		.reconfig_to_pll   (analyzer_pll_reconfig_reconfig_to_pll_reconfig_to_pll), //   reconfig_to_pll.reconfig_to_pll
		.reconfig_from_pll (analyzer_pll_reconfig_from_pll_reconfig_from_pll)       // reconfig_from_pll.reconfig_from_pll
	);

	altera_pll_reconfig_top #(
		.device_family       ("Cyclone V"),
		.ENABLE_MIF          (0),
		.MIF_FILE_NAME       (""),
		.ENABLE_BYTEENABLE   (0),
		.BYTEENABLE_WIDTH    (4),
		.RECONFIG_ADDR_WIDTH (6),
		.RECONFIG_DATA_WIDTH (32),
		.reconf_width        (64),
		.WAIT_FOR_LOCK       (1)
	) analyzer_pll_reconfig (
		.mgmt_clk          (clk_clk),                                                               //          mgmt_clk.clk
		.mgmt_reset        (rst_controller_003_reset_out_reset),                                    //        mgmt_reset.reset
		.mgmt_waitrequest  (mm_interconnect_1_analyzer_pll_reconfig_mgmt_avalon_slave_waitrequest), // mgmt_avalon_slave.waitrequest
		.mgmt_read         (mm_interconnect_1_analyzer_pll_reconfig_mgmt_avalon_slave_read),        //                  .read
		.mgmt_write        (mm_interconnect_1_analyzer_pll_reconfig_mgmt_avalon_slave_write),       //                  .write
		.mgmt_readdata     (mm_interconnect_1_analyzer_pll_reconfig_mgmt_avalon_slave_readdata),    //                  .readdata
		.mgmt_address      (mm_interconnect_1_analyzer_pll_reconfig_mgmt_avalon_slave_address),     //                  .address
		.mgmt_writedata    (mm_interconnect_1_analyzer_pll_reconfig_mgmt_avalon_slave_writedata),   //                  .writedata
		.reconfig_to_pll   (analyzer_pll_reconfig_reconfig_to_pll_reconfig_to_pll),                 //   reconfig_to_pll.reconfig_to_pll
		.reconfig_from_pll (analyzer_pll_reconfig_from_pll_reconfig_from_pll),                      // reconfig_from_pll.reconfig_from_pll
		.mgmt_byteenable   (4'b0000)                                                                //       (terminated)
	);

	soc_system_v5_aux_cnt_out aux_cnt_out (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_003_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_1_aux_cnt_out_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_aux_cnt_out_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_aux_cnt_out_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_aux_cnt_out_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_aux_cnt_out_s1_readdata),   //                    .readdata
		.out_port   (aux_cnt_out_export)                           // external_connection.export
	);

	soc_system_v5_ctrl_in ctrl_in (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_003_reset_out_reset),   //               reset.reset_n
		.address  (mm_interconnect_1_ctrl_in_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_ctrl_in_s1_readdata), //                    .readdata
		.in_port  (ctrl_in_export)                         // external_connection.export
	);

	soc_system_v5_aux_cnt_out ctrl_out (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_003_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_1_ctrl_out_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_ctrl_out_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_ctrl_out_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_ctrl_out_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_ctrl_out_s1_readdata),   //                    .readdata
		.out_port   (ctrl_out_export)                           // external_connection.export
	);

	soc_system_v5_dac_grad dac_grad (
		.clk           (clk_clk),                                                //              clk.clk
		.reset_n       (~rst_controller_003_reset_out_reset),                    //            reset.reset_n
		.data_from_cpu (mm_interconnect_1_dac_grad_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_1_dac_grad_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_1_dac_grad_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_1_dac_grad_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_1_dac_grad_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_1_dac_grad_spi_control_port_write),     //                 .write_n
		.irq           (irq_mapper_001_receiver2_irq),                           //              irq.irq
		.MISO          (dac_grad_MISO),                                          //         external.export
		.MOSI          (dac_grad_MOSI),                                          //                 .export
		.SCLK          (dac_grad_SCLK),                                          //                 .export
		.SS_n          (dac_grad_SS_n)                                           //                 .export
	);

	altera_avalon_dc_fifo #(
		.SYMBOLS_PER_BEAT   (1),
		.BITS_PER_SYMBOL    (32),
		.FIFO_DEPTH         (32768),
		.CHANNEL_WIDTH      (0),
		.ERROR_WIDTH        (0),
		.USE_PACKETS        (0),
		.USE_IN_FILL_LEVEL  (0),
		.USE_OUT_FILL_LEVEL (0),
		.WR_SYNC_DEPTH      (3),
		.RD_SYNC_DEPTH      (3)
	) dconv_fifo_dc (
		.in_clk            (fifo_clk_bridge_in_clk),               //        in_clk.clk
		.in_reset_n        (~rst_controller_reset_out_reset),      //  in_clk_reset.reset_n
		.out_clk           (clk_clk),                              //       out_clk.clk
		.out_reset_n       (~rst_controller_001_reset_out_reset),  // out_clk_reset.reset_n
		.in_data           (dconv_fifo_in_data),                   //            in.data
		.in_valid          (dconv_fifo_in_valid),                  //              .valid
		.in_ready          (dconv_fifo_in_ready),                  //              .ready
		.out_data          (dconv_fifo_dc_out_data),               //           out.data
		.out_valid         (dconv_fifo_dc_out_valid),              //              .valid
		.out_ready         (dconv_fifo_dc_out_ready),              //              .ready
		.in_csr_address    (1'b0),                                 //   (terminated)
		.in_csr_read       (1'b0),                                 //   (terminated)
		.in_csr_write      (1'b0),                                 //   (terminated)
		.in_csr_readdata   (),                                     //   (terminated)
		.in_csr_writedata  (32'b00000000000000000000000000000000), //   (terminated)
		.out_csr_address   (1'b0),                                 //   (terminated)
		.out_csr_read      (1'b0),                                 //   (terminated)
		.out_csr_write     (1'b0),                                 //   (terminated)
		.out_csr_readdata  (),                                     //   (terminated)
		.out_csr_writedata (32'b00000000000000000000000000000000), //   (terminated)
		.in_startofpacket  (1'b0),                                 //   (terminated)
		.in_endofpacket    (1'b0),                                 //   (terminated)
		.out_startofpacket (),                                     //   (terminated)
		.out_endofpacket   (),                                     //   (terminated)
		.in_empty          (1'b0),                                 //   (terminated)
		.out_empty         (),                                     //   (terminated)
		.in_error          (1'b0),                                 //   (terminated)
		.out_error         (),                                     //   (terminated)
		.in_channel        (1'b0),                                 //   (terminated)
		.out_channel       (),                                     //   (terminated)
		.space_avail_data  ()                                      //   (terminated)
	);

	altera_avalon_dc_fifo #(
		.SYMBOLS_PER_BEAT   (1),
		.BITS_PER_SYMBOL    (32),
		.FIFO_DEPTH         (32768),
		.CHANNEL_WIDTH      (0),
		.ERROR_WIDTH        (0),
		.USE_PACKETS        (0),
		.USE_IN_FILL_LEVEL  (0),
		.USE_OUT_FILL_LEVEL (0),
		.WR_SYNC_DEPTH      (3),
		.RD_SYNC_DEPTH      (3)
	) dconv_fifo_dc_q (
		.in_clk            (fifo_clk_bridge_in_clk),               //        in_clk.clk
		.in_reset_n        (~rst_controller_reset_out_reset),      //  in_clk_reset.reset_n
		.out_clk           (clk_clk),                              //       out_clk.clk
		.out_reset_n       (~rst_controller_001_reset_out_reset),  // out_clk_reset.reset_n
		.in_data           (dconv_fifo_q_in_data),                 //            in.data
		.in_valid          (dconv_fifo_q_in_valid),                //              .valid
		.in_ready          (dconv_fifo_q_in_ready),                //              .ready
		.out_data          (dconv_fifo_dc_q_out_data),             //           out.data
		.out_valid         (dconv_fifo_dc_q_out_valid),            //              .valid
		.out_ready         (dconv_fifo_dc_q_out_ready),            //              .ready
		.in_csr_address    (1'b0),                                 //   (terminated)
		.in_csr_read       (1'b0),                                 //   (terminated)
		.in_csr_write      (1'b0),                                 //   (terminated)
		.in_csr_readdata   (),                                     //   (terminated)
		.in_csr_writedata  (32'b00000000000000000000000000000000), //   (terminated)
		.out_csr_address   (1'b0),                                 //   (terminated)
		.out_csr_read      (1'b0),                                 //   (terminated)
		.out_csr_write     (1'b0),                                 //   (terminated)
		.out_csr_readdata  (),                                     //   (terminated)
		.out_csr_writedata (32'b00000000000000000000000000000000), //   (terminated)
		.in_startofpacket  (1'b0),                                 //   (terminated)
		.in_endofpacket    (1'b0),                                 //   (terminated)
		.out_startofpacket (),                                     //   (terminated)
		.out_endofpacket   (),                                     //   (terminated)
		.in_empty          (1'b0),                                 //   (terminated)
		.out_empty         (),                                     //   (terminated)
		.in_error          (1'b0),                                 //   (terminated)
		.out_error         (),                                     //   (terminated)
		.in_channel        (1'b0),                                 //   (terminated)
		.out_channel       (),                                     //   (terminated)
		.space_avail_data  ()                                      //   (terminated)
	);

	soc_system_v5_dconv_fifo_mem dconv_fifo_mem (
		.wrclock                         (clk_clk),                                           //   clk_in.clk
		.reset_n                         (~rst_controller_001_reset_out_reset),               // reset_in.reset_n
		.avalonst_sink_valid             (avalon_st_adapter_001_out_0_valid),                 //       in.valid
		.avalonst_sink_data              (avalon_st_adapter_001_out_0_data),                  //         .data
		.avalonst_sink_ready             (avalon_st_adapter_001_out_0_ready),                 //         .ready
		.avalonmm_read_slave_readdata    (mm_interconnect_1_dconv_fifo_mem_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read        (mm_interconnect_1_dconv_fifo_mem_out_read),         //         .read
		.avalonmm_read_slave_address     (mm_interconnect_1_dconv_fifo_mem_out_address),      //         .address
		.avalonmm_read_slave_waitrequest (mm_interconnect_1_dconv_fifo_mem_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address     (mm_interconnect_1_dconv_fifo_mem_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read        (mm_interconnect_1_dconv_fifo_mem_in_csr_read),      //         .read
		.wrclk_control_slave_writedata   (mm_interconnect_1_dconv_fifo_mem_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write       (mm_interconnect_1_dconv_fifo_mem_in_csr_write),     //         .write
		.wrclk_control_slave_readdata    (mm_interconnect_1_dconv_fifo_mem_in_csr_readdata)   //         .readdata
	);

	soc_system_v5_dconv_fifo_mem dconv_fifo_mem_q (
		.wrclock                         (clk_clk),                                             //   clk_in.clk
		.reset_n                         (~rst_controller_001_reset_out_reset),                 // reset_in.reset_n
		.avalonst_sink_valid             (avalon_st_adapter_002_out_0_valid),                   //       in.valid
		.avalonst_sink_data              (avalon_st_adapter_002_out_0_data),                    //         .data
		.avalonst_sink_ready             (avalon_st_adapter_002_out_0_ready),                   //         .ready
		.avalonmm_read_slave_readdata    (mm_interconnect_1_dconv_fifo_mem_q_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read        (mm_interconnect_1_dconv_fifo_mem_q_out_read),         //         .read
		.avalonmm_read_slave_address     (mm_interconnect_1_dconv_fifo_mem_q_out_address),      //         .address
		.avalonmm_read_slave_waitrequest (mm_interconnect_1_dconv_fifo_mem_q_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address     (mm_interconnect_1_dconv_fifo_mem_q_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read        (mm_interconnect_1_dconv_fifo_mem_q_in_csr_read),      //         .read
		.wrclk_control_slave_writedata   (mm_interconnect_1_dconv_fifo_mem_q_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write       (mm_interconnect_1_dconv_fifo_mem_q_in_csr_write),     //         .write
		.wrclk_control_slave_readdata    (mm_interconnect_1_dconv_fifo_mem_q_in_csr_readdata)   //         .readdata
	);

	soc_system_v5_dconv_fir dconv_fir (
		.clk              (fifo_clk_bridge_in_clk),                                    //                     clk.clk
		.reset_n          (~fifo_rst_reset),                                           //                     rst.reset_n
		.ast_sink_data    (dconv_fir_in_data),                                         //   avalon_streaming_sink.data
		.ast_sink_valid   (dconv_fir_in_valid),                                        //                        .valid
		.ast_sink_error   (dconv_fir_in_error),                                        //                        .error
		.ast_source_data  (dconv_fir_out_data),                                        // avalon_streaming_source.data
		.ast_source_valid (dconv_fir_out_valid),                                       //                        .valid
		.ast_source_error (dconv_fir_out_error),                                       //                        .error
		.coeff_in_clk     (clk_clk),                                                   //             coeff_clock.clk
		.coeff_in_areset  (~rst_controller_003_reset_out_reset),                       //             coeff_reset.reset_n
		.coeff_in_address (mm_interconnect_1_dconv_fir_avalon_mm_slave_address),       //         avalon_mm_slave.address
		.coeff_in_read    (mm_interconnect_1_dconv_fir_avalon_mm_slave_read),          //                        .read
		.coeff_out_valid  (mm_interconnect_1_dconv_fir_avalon_mm_slave_readdatavalid), //                        .readdatavalid
		.coeff_out_data   (mm_interconnect_1_dconv_fir_avalon_mm_slave_readdata),      //                        .readdata
		.coeff_in_we      (mm_interconnect_1_dconv_fir_avalon_mm_slave_write),         //                        .write
		.coeff_in_data    (mm_interconnect_1_dconv_fir_avalon_mm_slave_writedata)      //                        .writedata
	);

	soc_system_v5_dconv_fir dconv_fir_q (
		.clk              (fifo_clk_bridge_in_clk),                                      //                     clk.clk
		.reset_n          (~fifo_rst_reset),                                             //                     rst.reset_n
		.ast_sink_data    (dconv_fir_q_in_data),                                         //   avalon_streaming_sink.data
		.ast_sink_valid   (dconv_fir_q_in_valid),                                        //                        .valid
		.ast_sink_error   (dconv_fir_q_in_error),                                        //                        .error
		.ast_source_data  (dconv_fir_q_out_data),                                        // avalon_streaming_source.data
		.ast_source_valid (dconv_fir_q_out_valid),                                       //                        .valid
		.ast_source_error (dconv_fir_q_out_error),                                       //                        .error
		.coeff_in_clk     (clk_clk),                                                     //             coeff_clock.clk
		.coeff_in_areset  (~rst_controller_003_reset_out_reset),                         //             coeff_reset.reset_n
		.coeff_in_address (mm_interconnect_1_dconv_fir_q_avalon_mm_slave_address),       //         avalon_mm_slave.address
		.coeff_in_read    (mm_interconnect_1_dconv_fir_q_avalon_mm_slave_read),          //                        .read
		.coeff_out_valid  (mm_interconnect_1_dconv_fir_q_avalon_mm_slave_readdatavalid), //                        .readdatavalid
		.coeff_out_data   (mm_interconnect_1_dconv_fir_q_avalon_mm_slave_readdata),      //                        .readdata
		.coeff_in_we      (mm_interconnect_1_dconv_fir_q_avalon_mm_slave_write),         //                        .write
		.coeff_in_data    (mm_interconnect_1_dconv_fir_q_avalon_mm_slave_writedata)      //                        .writedata
	);

	soc_system_v5_dma_dconvi dma_dconvi (
		.clk                (clk_clk),                                                    //                clk.clk
		.system_reset_n     (~rst_controller_003_reset_out_reset),                        //              reset.reset_n
		.dma_ctl_address    (mm_interconnect_1_dma_dconvi_control_port_slave_address),    // control_port_slave.address
		.dma_ctl_chipselect (mm_interconnect_1_dma_dconvi_control_port_slave_chipselect), //                   .chipselect
		.dma_ctl_readdata   (mm_interconnect_1_dma_dconvi_control_port_slave_readdata),   //                   .readdata
		.dma_ctl_write_n    (~mm_interconnect_1_dma_dconvi_control_port_slave_write),     //                   .write_n
		.dma_ctl_writedata  (mm_interconnect_1_dma_dconvi_control_port_slave_writedata),  //                   .writedata
		.dma_ctl_irq        (irq_mapper_001_receiver5_irq),                               //                irq.irq
		.read_address       (dma_dconvi_read_master_address),                             //        read_master.address
		.read_chipselect    (dma_dconvi_read_master_chipselect),                          //                   .chipselect
		.read_read_n        (dma_dconvi_read_master_read),                                //                   .read_n
		.read_readdata      (dma_dconvi_read_master_readdata),                            //                   .readdata
		.read_readdatavalid (dma_dconvi_read_master_readdatavalid),                       //                   .readdatavalid
		.read_waitrequest   (dma_dconvi_read_master_waitrequest),                         //                   .waitrequest
		.write_address      (dma_dconvi_write_master_address),                            //       write_master.address
		.write_chipselect   (dma_dconvi_write_master_chipselect),                         //                   .chipselect
		.write_waitrequest  (dma_dconvi_write_master_waitrequest),                        //                   .waitrequest
		.write_write_n      (dma_dconvi_write_master_write),                              //                   .write_n
		.write_writedata    (dma_dconvi_write_master_writedata),                          //                   .writedata
		.write_byteenable   (dma_dconvi_write_master_byteenable)                          //                   .byteenable
	);

	soc_system_v5_dma_dconvq dma_dconvq (
		.clk                (clk_clk),                                                    //                clk.clk
		.system_reset_n     (~rst_controller_003_reset_out_reset),                        //              reset.reset_n
		.dma_ctl_address    (mm_interconnect_1_dma_dconvq_control_port_slave_address),    // control_port_slave.address
		.dma_ctl_chipselect (mm_interconnect_1_dma_dconvq_control_port_slave_chipselect), //                   .chipselect
		.dma_ctl_readdata   (mm_interconnect_1_dma_dconvq_control_port_slave_readdata),   //                   .readdata
		.dma_ctl_write_n    (~mm_interconnect_1_dma_dconvq_control_port_slave_write),     //                   .write_n
		.dma_ctl_writedata  (mm_interconnect_1_dma_dconvq_control_port_slave_writedata),  //                   .writedata
		.dma_ctl_irq        (irq_mapper_001_receiver6_irq),                               //                irq.irq
		.read_address       (dma_dconvq_read_master_address),                             //        read_master.address
		.read_chipselect    (dma_dconvq_read_master_chipselect),                          //                   .chipselect
		.read_read_n        (dma_dconvq_read_master_read),                                //                   .read_n
		.read_readdata      (dma_dconvq_read_master_readdata),                            //                   .readdata
		.read_readdatavalid (dma_dconvq_read_master_readdatavalid),                       //                   .readdatavalid
		.read_waitrequest   (dma_dconvq_read_master_waitrequest),                         //                   .waitrequest
		.write_address      (dma_dconvq_write_master_address),                            //       write_master.address
		.write_chipselect   (dma_dconvq_write_master_chipselect),                         //                   .chipselect
		.write_waitrequest  (dma_dconvq_write_master_waitrequest),                        //                   .waitrequest
		.write_write_n      (dma_dconvq_write_master_write),                              //                   .write_n
		.write_writedata    (dma_dconvq_write_master_writedata),                          //                   .writedata
		.write_byteenable   (dma_dconvq_write_master_byteenable)                          //                   .byteenable
	);

	soc_system_v5_dma_dummy dma_dummy (
		.clk                (clk_clk),                                                   //                clk.clk
		.system_reset_n     (~rst_controller_003_reset_out_reset),                       //              reset.reset_n
		.dma_ctl_address    (mm_interconnect_1_dma_dummy_control_port_slave_address),    // control_port_slave.address
		.dma_ctl_chipselect (mm_interconnect_1_dma_dummy_control_port_slave_chipselect), //                   .chipselect
		.dma_ctl_readdata   (mm_interconnect_1_dma_dummy_control_port_slave_readdata),   //                   .readdata
		.dma_ctl_write_n    (~mm_interconnect_1_dma_dummy_control_port_slave_write),     //                   .write_n
		.dma_ctl_writedata  (mm_interconnect_1_dma_dummy_control_port_slave_writedata),  //                   .writedata
		.dma_ctl_irq        (),                                                          //                irq.irq
		.read_address       (dma_dummy_read_master_address),                             //        read_master.address
		.read_chipselect    (dma_dummy_read_master_chipselect),                          //                   .chipselect
		.read_read_n        (dma_dummy_read_master_read),                                //                   .read_n
		.read_readdata      (dma_dummy_read_master_readdata),                            //                   .readdata
		.read_readdatavalid (dma_dummy_read_master_readdatavalid),                       //                   .readdatavalid
		.read_waitrequest   (dma_dummy_read_master_waitrequest),                         //                   .waitrequest
		.write_address      (dma_dummy_write_master_address),                            //       write_master.address
		.write_chipselect   (dma_dummy_write_master_chipselect),                         //                   .chipselect
		.write_waitrequest  (dma_dummy_write_master_waitrequest),                        //                   .waitrequest
		.write_write_n      (dma_dummy_write_master_write),                              //                   .write_n
		.write_writedata    (dma_dummy_write_master_writedata),                          //                   .writedata
		.write_byteenable   (dma_dummy_write_master_byteenable)                          //                   .byteenable
	);

	soc_system_v5_dma_fifo dma_fifo (
		.clk                (clk_clk),                                                  //                clk.clk
		.system_reset_n     (~rst_controller_003_reset_out_reset),                      //              reset.reset_n
		.dma_ctl_address    (mm_interconnect_1_dma_fifo_control_port_slave_address),    // control_port_slave.address
		.dma_ctl_chipselect (mm_interconnect_1_dma_fifo_control_port_slave_chipselect), //                   .chipselect
		.dma_ctl_readdata   (mm_interconnect_1_dma_fifo_control_port_slave_readdata),   //                   .readdata
		.dma_ctl_write_n    (~mm_interconnect_1_dma_fifo_control_port_slave_write),     //                   .write_n
		.dma_ctl_writedata  (mm_interconnect_1_dma_fifo_control_port_slave_writedata),  //                   .writedata
		.dma_ctl_irq        (irq_mapper_001_receiver3_irq),                             //                irq.irq
		.read_address       (dma_fifo_read_master_address),                             //        read_master.address
		.read_chipselect    (dma_fifo_read_master_chipselect),                          //                   .chipselect
		.read_read_n        (dma_fifo_read_master_read),                                //                   .read_n
		.read_readdata      (dma_fifo_read_master_readdata),                            //                   .readdata
		.read_readdatavalid (dma_fifo_read_master_readdatavalid),                       //                   .readdatavalid
		.read_waitrequest   (dma_fifo_read_master_waitrequest),                         //                   .waitrequest
		.write_address      (dma_fifo_write_master_address),                            //       write_master.address
		.write_chipselect   (dma_fifo_write_master_chipselect),                         //                   .chipselect
		.write_waitrequest  (dma_fifo_write_master_waitrequest),                        //                   .waitrequest
		.write_write_n      (dma_fifo_write_master_write),                              //                   .write_n
		.write_writedata    (dma_fifo_write_master_writedata),                          //                   .writedata
		.write_byteenable   (dma_fifo_write_master_byteenable)                          //                   .byteenable
	);

	soc_system_v5_fifo_dummy fifo_dummy (
		.wrclock                          (clk_clk),                                       //   clk_in.clk
		.reset_n                          (~rst_controller_003_reset_out_reset),           // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_1_fifo_dummy_in_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_1_fifo_dummy_in_write),         //         .write
		.avalonmm_write_slave_waitrequest (mm_interconnect_1_fifo_dummy_in_waitrequest),   //         .waitrequest
		.avalonmm_read_slave_readdata     (mm_interconnect_1_fifo_dummy_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (mm_interconnect_1_fifo_dummy_out_read),         //         .read
		.avalonmm_read_slave_waitrequest  (mm_interconnect_1_fifo_dummy_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address      (mm_interconnect_1_fifo_dummy_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_1_fifo_dummy_in_csr_read),      //         .read
		.wrclk_control_slave_writedata    (mm_interconnect_1_fifo_dummy_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write        (mm_interconnect_1_fifo_dummy_in_csr_write),     //         .write
		.wrclk_control_slave_readdata     (mm_interconnect_1_fifo_dummy_in_csr_readdata)   //         .readdata
	);

	soc_system_v5_fifo_dummy64_in fifo_dummy64_in (
		.wrclock                          (clk_clk),                                            //   clk_in.clk
		.reset_n                          (~rst_controller_003_reset_out_reset),                // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_1_fifo_dummy64_in_in_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_1_fifo_dummy64_in_in_write),         //         .write
		.avalonmm_write_slave_address     (mm_interconnect_1_fifo_dummy64_in_in_address),       //         .address
		.avalonmm_write_slave_waitrequest (mm_interconnect_1_fifo_dummy64_in_in_waitrequest),   //         .waitrequest
		.avalonst_source_valid            (fifo_dummy64_in_out_valid),                          //      out.valid
		.avalonst_source_data             (fifo_dummy64_in_out_data),                           //         .data
		.avalonst_source_ready            (fifo_dummy64_in_out_ready),                          //         .ready
		.wrclk_control_slave_address      (mm_interconnect_1_fifo_dummy64_in_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_1_fifo_dummy64_in_in_csr_read),      //         .read
		.wrclk_control_slave_writedata    (mm_interconnect_1_fifo_dummy64_in_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write        (mm_interconnect_1_fifo_dummy64_in_in_csr_write),     //         .write
		.wrclk_control_slave_readdata     (mm_interconnect_1_fifo_dummy64_in_in_csr_readdata)   //         .readdata
	);

	soc_system_v5_fifo_dummy64_out fifo_dummy64_out (
		.wrclock                         (clk_clk),                                             //   clk_in.clk
		.reset_n                         (~rst_controller_003_reset_out_reset),                 // reset_in.reset_n
		.avalonst_sink_valid             (fifo_dummy64_in_out_valid),                           //       in.valid
		.avalonst_sink_data              (fifo_dummy64_in_out_data),                            //         .data
		.avalonst_sink_ready             (fifo_dummy64_in_out_ready),                           //         .ready
		.avalonmm_read_slave_readdata    (mm_interconnect_1_fifo_dummy64_out_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read        (mm_interconnect_1_fifo_dummy64_out_out_read),         //         .read
		.avalonmm_read_slave_address     (mm_interconnect_1_fifo_dummy64_out_out_address),      //         .address
		.avalonmm_read_slave_waitrequest (mm_interconnect_1_fifo_dummy64_out_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address     (mm_interconnect_1_fifo_dummy64_out_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read        (mm_interconnect_1_fifo_dummy64_out_in_csr_read),      //         .read
		.wrclk_control_slave_writedata   (mm_interconnect_1_fifo_dummy64_out_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write       (mm_interconnect_1_fifo_dummy64_out_in_csr_write),     //         .write
		.wrclk_control_slave_readdata    (mm_interconnect_1_fifo_dummy64_out_in_csr_readdata)   //         .readdata
	);

	soc_system_v5_gp_pll gp_pll (
		.refclk   (clk_clk),               //  refclk.clk
		.rst      (~reset_reset_n),        //   reset.reset
		.outclk_0 (gp_pll_outclk0_clk),    // outclk0.clk
		.outclk_1 (pll_vga_clk65_clk),     // outclk1.clk
		.outclk_2 (),                      // outclk2.clk
		.outclk_3 (sdram_clk_clk),         // outclk3.clk
		.locked   (pll_vga_locked_export)  //  locked.export
	);

	soc_system_v5_hps_0 #(
		.F2S_Width (3),
		.S2F_Width (3)
	) hps_0 (
		.mem_a                    (memory_mem_a),                                  //            memory.mem_a
		.mem_ba                   (memory_mem_ba),                                 //                  .mem_ba
		.mem_ck                   (memory_mem_ck),                                 //                  .mem_ck
		.mem_ck_n                 (memory_mem_ck_n),                               //                  .mem_ck_n
		.mem_cke                  (memory_mem_cke),                                //                  .mem_cke
		.mem_cs_n                 (memory_mem_cs_n),                               //                  .mem_cs_n
		.mem_ras_n                (memory_mem_ras_n),                              //                  .mem_ras_n
		.mem_cas_n                (memory_mem_cas_n),                              //                  .mem_cas_n
		.mem_we_n                 (memory_mem_we_n),                               //                  .mem_we_n
		.mem_reset_n              (memory_mem_reset_n),                            //                  .mem_reset_n
		.mem_dq                   (memory_mem_dq),                                 //                  .mem_dq
		.mem_dqs                  (memory_mem_dqs),                                //                  .mem_dqs
		.mem_dqs_n                (memory_mem_dqs_n),                              //                  .mem_dqs_n
		.mem_odt                  (memory_mem_odt),                                //                  .mem_odt
		.mem_dm                   (memory_mem_dm),                                 //                  .mem_dm
		.oct_rzqin                (memory_oct_rzqin),                              //                  .oct_rzqin
		.hps_io_emac1_inst_TX_CLK (hps_0_hps_io_hps_io_emac1_inst_TX_CLK),         //            hps_io.hps_io_emac1_inst_TX_CLK
		.hps_io_emac1_inst_TXD0   (hps_0_hps_io_hps_io_emac1_inst_TXD0),           //                  .hps_io_emac1_inst_TXD0
		.hps_io_emac1_inst_TXD1   (hps_0_hps_io_hps_io_emac1_inst_TXD1),           //                  .hps_io_emac1_inst_TXD1
		.hps_io_emac1_inst_TXD2   (hps_0_hps_io_hps_io_emac1_inst_TXD2),           //                  .hps_io_emac1_inst_TXD2
		.hps_io_emac1_inst_TXD3   (hps_0_hps_io_hps_io_emac1_inst_TXD3),           //                  .hps_io_emac1_inst_TXD3
		.hps_io_emac1_inst_RXD0   (hps_0_hps_io_hps_io_emac1_inst_RXD0),           //                  .hps_io_emac1_inst_RXD0
		.hps_io_emac1_inst_MDIO   (hps_0_hps_io_hps_io_emac1_inst_MDIO),           //                  .hps_io_emac1_inst_MDIO
		.hps_io_emac1_inst_MDC    (hps_0_hps_io_hps_io_emac1_inst_MDC),            //                  .hps_io_emac1_inst_MDC
		.hps_io_emac1_inst_RX_CTL (hps_0_hps_io_hps_io_emac1_inst_RX_CTL),         //                  .hps_io_emac1_inst_RX_CTL
		.hps_io_emac1_inst_TX_CTL (hps_0_hps_io_hps_io_emac1_inst_TX_CTL),         //                  .hps_io_emac1_inst_TX_CTL
		.hps_io_emac1_inst_RX_CLK (hps_0_hps_io_hps_io_emac1_inst_RX_CLK),         //                  .hps_io_emac1_inst_RX_CLK
		.hps_io_emac1_inst_RXD1   (hps_0_hps_io_hps_io_emac1_inst_RXD1),           //                  .hps_io_emac1_inst_RXD1
		.hps_io_emac1_inst_RXD2   (hps_0_hps_io_hps_io_emac1_inst_RXD2),           //                  .hps_io_emac1_inst_RXD2
		.hps_io_emac1_inst_RXD3   (hps_0_hps_io_hps_io_emac1_inst_RXD3),           //                  .hps_io_emac1_inst_RXD3
		.hps_io_qspi_inst_IO0     (hps_0_hps_io_hps_io_qspi_inst_IO0),             //                  .hps_io_qspi_inst_IO0
		.hps_io_qspi_inst_IO1     (hps_0_hps_io_hps_io_qspi_inst_IO1),             //                  .hps_io_qspi_inst_IO1
		.hps_io_qspi_inst_IO2     (hps_0_hps_io_hps_io_qspi_inst_IO2),             //                  .hps_io_qspi_inst_IO2
		.hps_io_qspi_inst_IO3     (hps_0_hps_io_hps_io_qspi_inst_IO3),             //                  .hps_io_qspi_inst_IO3
		.hps_io_qspi_inst_SS0     (hps_0_hps_io_hps_io_qspi_inst_SS0),             //                  .hps_io_qspi_inst_SS0
		.hps_io_qspi_inst_CLK     (hps_0_hps_io_hps_io_qspi_inst_CLK),             //                  .hps_io_qspi_inst_CLK
		.hps_io_sdio_inst_CMD     (hps_0_hps_io_hps_io_sdio_inst_CMD),             //                  .hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0      (hps_0_hps_io_hps_io_sdio_inst_D0),              //                  .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1      (hps_0_hps_io_hps_io_sdio_inst_D1),              //                  .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK     (hps_0_hps_io_hps_io_sdio_inst_CLK),             //                  .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2      (hps_0_hps_io_hps_io_sdio_inst_D2),              //                  .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3      (hps_0_hps_io_hps_io_sdio_inst_D3),              //                  .hps_io_sdio_inst_D3
		.hps_io_usb1_inst_D0      (hps_0_hps_io_hps_io_usb1_inst_D0),              //                  .hps_io_usb1_inst_D0
		.hps_io_usb1_inst_D1      (hps_0_hps_io_hps_io_usb1_inst_D1),              //                  .hps_io_usb1_inst_D1
		.hps_io_usb1_inst_D2      (hps_0_hps_io_hps_io_usb1_inst_D2),              //                  .hps_io_usb1_inst_D2
		.hps_io_usb1_inst_D3      (hps_0_hps_io_hps_io_usb1_inst_D3),              //                  .hps_io_usb1_inst_D3
		.hps_io_usb1_inst_D4      (hps_0_hps_io_hps_io_usb1_inst_D4),              //                  .hps_io_usb1_inst_D4
		.hps_io_usb1_inst_D5      (hps_0_hps_io_hps_io_usb1_inst_D5),              //                  .hps_io_usb1_inst_D5
		.hps_io_usb1_inst_D6      (hps_0_hps_io_hps_io_usb1_inst_D6),              //                  .hps_io_usb1_inst_D6
		.hps_io_usb1_inst_D7      (hps_0_hps_io_hps_io_usb1_inst_D7),              //                  .hps_io_usb1_inst_D7
		.hps_io_usb1_inst_CLK     (hps_0_hps_io_hps_io_usb1_inst_CLK),             //                  .hps_io_usb1_inst_CLK
		.hps_io_usb1_inst_STP     (hps_0_hps_io_hps_io_usb1_inst_STP),             //                  .hps_io_usb1_inst_STP
		.hps_io_usb1_inst_DIR     (hps_0_hps_io_hps_io_usb1_inst_DIR),             //                  .hps_io_usb1_inst_DIR
		.hps_io_usb1_inst_NXT     (hps_0_hps_io_hps_io_usb1_inst_NXT),             //                  .hps_io_usb1_inst_NXT
		.hps_io_spim1_inst_CLK    (hps_0_hps_io_hps_io_spim1_inst_CLK),            //                  .hps_io_spim1_inst_CLK
		.hps_io_spim1_inst_MOSI   (hps_0_hps_io_hps_io_spim1_inst_MOSI),           //                  .hps_io_spim1_inst_MOSI
		.hps_io_spim1_inst_MISO   (hps_0_hps_io_hps_io_spim1_inst_MISO),           //                  .hps_io_spim1_inst_MISO
		.hps_io_spim1_inst_SS0    (hps_0_hps_io_hps_io_spim1_inst_SS0),            //                  .hps_io_spim1_inst_SS0
		.hps_io_uart0_inst_RX     (hps_0_hps_io_hps_io_uart0_inst_RX),             //                  .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX     (hps_0_hps_io_hps_io_uart0_inst_TX),             //                  .hps_io_uart0_inst_TX
		.hps_io_i2c0_inst_SDA     (hps_0_hps_io_hps_io_i2c0_inst_SDA),             //                  .hps_io_i2c0_inst_SDA
		.hps_io_i2c0_inst_SCL     (hps_0_hps_io_hps_io_i2c0_inst_SCL),             //                  .hps_io_i2c0_inst_SCL
		.hps_io_i2c1_inst_SDA     (hps_0_hps_io_hps_io_i2c1_inst_SDA),             //                  .hps_io_i2c1_inst_SDA
		.hps_io_i2c1_inst_SCL     (hps_0_hps_io_hps_io_i2c1_inst_SCL),             //                  .hps_io_i2c1_inst_SCL
		.hps_io_gpio_inst_GPIO09  (hps_0_hps_io_hps_io_gpio_inst_GPIO09),          //                  .hps_io_gpio_inst_GPIO09
		.hps_io_gpio_inst_GPIO35  (hps_0_hps_io_hps_io_gpio_inst_GPIO35),          //                  .hps_io_gpio_inst_GPIO35
		.hps_io_gpio_inst_GPIO40  (hps_0_hps_io_hps_io_gpio_inst_GPIO40),          //                  .hps_io_gpio_inst_GPIO40
		.hps_io_gpio_inst_GPIO48  (hps_0_hps_io_hps_io_gpio_inst_GPIO48),          //                  .hps_io_gpio_inst_GPIO48
		.hps_io_gpio_inst_GPIO53  (hps_0_hps_io_hps_io_gpio_inst_GPIO53),          //                  .hps_io_gpio_inst_GPIO53
		.hps_io_gpio_inst_GPIO54  (hps_0_hps_io_hps_io_gpio_inst_GPIO54),          //                  .hps_io_gpio_inst_GPIO54
		.hps_io_gpio_inst_GPIO61  (hps_0_hps_io_hps_io_gpio_inst_GPIO61),          //                  .hps_io_gpio_inst_GPIO61
		.h2f_rst_n                (hps_0_h2f_reset_reset_n),                       //         h2f_reset.reset_n
		.h2f_axi_clk              (clk_clk),                                       //     h2f_axi_clock.clk
		.h2f_AWID                 (hps_0_h2f_axi_master_awid),                     //    h2f_axi_master.awid
		.h2f_AWADDR               (hps_0_h2f_axi_master_awaddr),                   //                  .awaddr
		.h2f_AWLEN                (hps_0_h2f_axi_master_awlen),                    //                  .awlen
		.h2f_AWSIZE               (hps_0_h2f_axi_master_awsize),                   //                  .awsize
		.h2f_AWBURST              (hps_0_h2f_axi_master_awburst),                  //                  .awburst
		.h2f_AWLOCK               (hps_0_h2f_axi_master_awlock),                   //                  .awlock
		.h2f_AWCACHE              (hps_0_h2f_axi_master_awcache),                  //                  .awcache
		.h2f_AWPROT               (hps_0_h2f_axi_master_awprot),                   //                  .awprot
		.h2f_AWVALID              (hps_0_h2f_axi_master_awvalid),                  //                  .awvalid
		.h2f_AWREADY              (hps_0_h2f_axi_master_awready),                  //                  .awready
		.h2f_WID                  (hps_0_h2f_axi_master_wid),                      //                  .wid
		.h2f_WDATA                (hps_0_h2f_axi_master_wdata),                    //                  .wdata
		.h2f_WSTRB                (hps_0_h2f_axi_master_wstrb),                    //                  .wstrb
		.h2f_WLAST                (hps_0_h2f_axi_master_wlast),                    //                  .wlast
		.h2f_WVALID               (hps_0_h2f_axi_master_wvalid),                   //                  .wvalid
		.h2f_WREADY               (hps_0_h2f_axi_master_wready),                   //                  .wready
		.h2f_BID                  (hps_0_h2f_axi_master_bid),                      //                  .bid
		.h2f_BRESP                (hps_0_h2f_axi_master_bresp),                    //                  .bresp
		.h2f_BVALID               (hps_0_h2f_axi_master_bvalid),                   //                  .bvalid
		.h2f_BREADY               (hps_0_h2f_axi_master_bready),                   //                  .bready
		.h2f_ARID                 (hps_0_h2f_axi_master_arid),                     //                  .arid
		.h2f_ARADDR               (hps_0_h2f_axi_master_araddr),                   //                  .araddr
		.h2f_ARLEN                (hps_0_h2f_axi_master_arlen),                    //                  .arlen
		.h2f_ARSIZE               (hps_0_h2f_axi_master_arsize),                   //                  .arsize
		.h2f_ARBURST              (hps_0_h2f_axi_master_arburst),                  //                  .arburst
		.h2f_ARLOCK               (hps_0_h2f_axi_master_arlock),                   //                  .arlock
		.h2f_ARCACHE              (hps_0_h2f_axi_master_arcache),                  //                  .arcache
		.h2f_ARPROT               (hps_0_h2f_axi_master_arprot),                   //                  .arprot
		.h2f_ARVALID              (hps_0_h2f_axi_master_arvalid),                  //                  .arvalid
		.h2f_ARREADY              (hps_0_h2f_axi_master_arready),                  //                  .arready
		.h2f_RID                  (hps_0_h2f_axi_master_rid),                      //                  .rid
		.h2f_RDATA                (hps_0_h2f_axi_master_rdata),                    //                  .rdata
		.h2f_RRESP                (hps_0_h2f_axi_master_rresp),                    //                  .rresp
		.h2f_RLAST                (hps_0_h2f_axi_master_rlast),                    //                  .rlast
		.h2f_RVALID               (hps_0_h2f_axi_master_rvalid),                   //                  .rvalid
		.h2f_RREADY               (hps_0_h2f_axi_master_rready),                   //                  .rready
		.f2h_axi_clk              (clk_clk),                                       //     f2h_axi_clock.clk
		.f2h_AWID                 (mm_interconnect_0_hps_0_f2h_axi_slave_awid),    //     f2h_axi_slave.awid
		.f2h_AWADDR               (mm_interconnect_0_hps_0_f2h_axi_slave_awaddr),  //                  .awaddr
		.f2h_AWLEN                (mm_interconnect_0_hps_0_f2h_axi_slave_awlen),   //                  .awlen
		.f2h_AWSIZE               (mm_interconnect_0_hps_0_f2h_axi_slave_awsize),  //                  .awsize
		.f2h_AWBURST              (mm_interconnect_0_hps_0_f2h_axi_slave_awburst), //                  .awburst
		.f2h_AWLOCK               (mm_interconnect_0_hps_0_f2h_axi_slave_awlock),  //                  .awlock
		.f2h_AWCACHE              (mm_interconnect_0_hps_0_f2h_axi_slave_awcache), //                  .awcache
		.f2h_AWPROT               (mm_interconnect_0_hps_0_f2h_axi_slave_awprot),  //                  .awprot
		.f2h_AWVALID              (mm_interconnect_0_hps_0_f2h_axi_slave_awvalid), //                  .awvalid
		.f2h_AWREADY              (mm_interconnect_0_hps_0_f2h_axi_slave_awready), //                  .awready
		.f2h_AWUSER               (mm_interconnect_0_hps_0_f2h_axi_slave_awuser),  //                  .awuser
		.f2h_WID                  (mm_interconnect_0_hps_0_f2h_axi_slave_wid),     //                  .wid
		.f2h_WDATA                (mm_interconnect_0_hps_0_f2h_axi_slave_wdata),   //                  .wdata
		.f2h_WSTRB                (mm_interconnect_0_hps_0_f2h_axi_slave_wstrb),   //                  .wstrb
		.f2h_WLAST                (mm_interconnect_0_hps_0_f2h_axi_slave_wlast),   //                  .wlast
		.f2h_WVALID               (mm_interconnect_0_hps_0_f2h_axi_slave_wvalid),  //                  .wvalid
		.f2h_WREADY               (mm_interconnect_0_hps_0_f2h_axi_slave_wready),  //                  .wready
		.f2h_BID                  (mm_interconnect_0_hps_0_f2h_axi_slave_bid),     //                  .bid
		.f2h_BRESP                (mm_interconnect_0_hps_0_f2h_axi_slave_bresp),   //                  .bresp
		.f2h_BVALID               (mm_interconnect_0_hps_0_f2h_axi_slave_bvalid),  //                  .bvalid
		.f2h_BREADY               (mm_interconnect_0_hps_0_f2h_axi_slave_bready),  //                  .bready
		.f2h_ARID                 (mm_interconnect_0_hps_0_f2h_axi_slave_arid),    //                  .arid
		.f2h_ARADDR               (mm_interconnect_0_hps_0_f2h_axi_slave_araddr),  //                  .araddr
		.f2h_ARLEN                (mm_interconnect_0_hps_0_f2h_axi_slave_arlen),   //                  .arlen
		.f2h_ARSIZE               (mm_interconnect_0_hps_0_f2h_axi_slave_arsize),  //                  .arsize
		.f2h_ARBURST              (mm_interconnect_0_hps_0_f2h_axi_slave_arburst), //                  .arburst
		.f2h_ARLOCK               (mm_interconnect_0_hps_0_f2h_axi_slave_arlock),  //                  .arlock
		.f2h_ARCACHE              (mm_interconnect_0_hps_0_f2h_axi_slave_arcache), //                  .arcache
		.f2h_ARPROT               (mm_interconnect_0_hps_0_f2h_axi_slave_arprot),  //                  .arprot
		.f2h_ARVALID              (mm_interconnect_0_hps_0_f2h_axi_slave_arvalid), //                  .arvalid
		.f2h_ARREADY              (mm_interconnect_0_hps_0_f2h_axi_slave_arready), //                  .arready
		.f2h_ARUSER               (mm_interconnect_0_hps_0_f2h_axi_slave_aruser),  //                  .aruser
		.f2h_RID                  (mm_interconnect_0_hps_0_f2h_axi_slave_rid),     //                  .rid
		.f2h_RDATA                (mm_interconnect_0_hps_0_f2h_axi_slave_rdata),   //                  .rdata
		.f2h_RRESP                (mm_interconnect_0_hps_0_f2h_axi_slave_rresp),   //                  .rresp
		.f2h_RLAST                (mm_interconnect_0_hps_0_f2h_axi_slave_rlast),   //                  .rlast
		.f2h_RVALID               (mm_interconnect_0_hps_0_f2h_axi_slave_rvalid),  //                  .rvalid
		.f2h_RREADY               (mm_interconnect_0_hps_0_f2h_axi_slave_rready),  //                  .rready
		.h2f_lw_axi_clk           (clk_clk),                                       //  h2f_lw_axi_clock.clk
		.h2f_lw_AWID              (hps_0_h2f_lw_axi_master_awid),                  // h2f_lw_axi_master.awid
		.h2f_lw_AWADDR            (hps_0_h2f_lw_axi_master_awaddr),                //                  .awaddr
		.h2f_lw_AWLEN             (hps_0_h2f_lw_axi_master_awlen),                 //                  .awlen
		.h2f_lw_AWSIZE            (hps_0_h2f_lw_axi_master_awsize),                //                  .awsize
		.h2f_lw_AWBURST           (hps_0_h2f_lw_axi_master_awburst),               //                  .awburst
		.h2f_lw_AWLOCK            (hps_0_h2f_lw_axi_master_awlock),                //                  .awlock
		.h2f_lw_AWCACHE           (hps_0_h2f_lw_axi_master_awcache),               //                  .awcache
		.h2f_lw_AWPROT            (hps_0_h2f_lw_axi_master_awprot),                //                  .awprot
		.h2f_lw_AWVALID           (hps_0_h2f_lw_axi_master_awvalid),               //                  .awvalid
		.h2f_lw_AWREADY           (hps_0_h2f_lw_axi_master_awready),               //                  .awready
		.h2f_lw_WID               (hps_0_h2f_lw_axi_master_wid),                   //                  .wid
		.h2f_lw_WDATA             (hps_0_h2f_lw_axi_master_wdata),                 //                  .wdata
		.h2f_lw_WSTRB             (hps_0_h2f_lw_axi_master_wstrb),                 //                  .wstrb
		.h2f_lw_WLAST             (hps_0_h2f_lw_axi_master_wlast),                 //                  .wlast
		.h2f_lw_WVALID            (hps_0_h2f_lw_axi_master_wvalid),                //                  .wvalid
		.h2f_lw_WREADY            (hps_0_h2f_lw_axi_master_wready),                //                  .wready
		.h2f_lw_BID               (hps_0_h2f_lw_axi_master_bid),                   //                  .bid
		.h2f_lw_BRESP             (hps_0_h2f_lw_axi_master_bresp),                 //                  .bresp
		.h2f_lw_BVALID            (hps_0_h2f_lw_axi_master_bvalid),                //                  .bvalid
		.h2f_lw_BREADY            (hps_0_h2f_lw_axi_master_bready),                //                  .bready
		.h2f_lw_ARID              (hps_0_h2f_lw_axi_master_arid),                  //                  .arid
		.h2f_lw_ARADDR            (hps_0_h2f_lw_axi_master_araddr),                //                  .araddr
		.h2f_lw_ARLEN             (hps_0_h2f_lw_axi_master_arlen),                 //                  .arlen
		.h2f_lw_ARSIZE            (hps_0_h2f_lw_axi_master_arsize),                //                  .arsize
		.h2f_lw_ARBURST           (hps_0_h2f_lw_axi_master_arburst),               //                  .arburst
		.h2f_lw_ARLOCK            (hps_0_h2f_lw_axi_master_arlock),                //                  .arlock
		.h2f_lw_ARCACHE           (hps_0_h2f_lw_axi_master_arcache),               //                  .arcache
		.h2f_lw_ARPROT            (hps_0_h2f_lw_axi_master_arprot),                //                  .arprot
		.h2f_lw_ARVALID           (hps_0_h2f_lw_axi_master_arvalid),               //                  .arvalid
		.h2f_lw_ARREADY           (hps_0_h2f_lw_axi_master_arready),               //                  .arready
		.h2f_lw_RID               (hps_0_h2f_lw_axi_master_rid),                   //                  .rid
		.h2f_lw_RDATA             (hps_0_h2f_lw_axi_master_rdata),                 //                  .rdata
		.h2f_lw_RRESP             (hps_0_h2f_lw_axi_master_rresp),                 //                  .rresp
		.h2f_lw_RLAST             (hps_0_h2f_lw_axi_master_rlast),                 //                  .rlast
		.h2f_lw_RVALID            (hps_0_h2f_lw_axi_master_rvalid),                //                  .rvalid
		.h2f_lw_RREADY            (hps_0_h2f_lw_axi_master_rready),                //                  .rready
		.f2h_irq_p0               (hps_0_f2h_irq0_irq),                            //          f2h_irq0.irq
		.f2h_irq_p1               (hps_0_f2h_irq1_irq)                             //          f2h_irq1.irq
	);

	altera_avalon_i2c #(
		.USE_AV_ST       (0),
		.FIFO_DEPTH      (32),
		.FIFO_DEPTH_LOG2 (5)
	) i2c_ext (
		.clk       (clk_clk),                                 //            clock.clk
		.rst_n     (~rst_controller_003_reset_out_reset),     //       reset_sink.reset_n
		.intr      (irq_mapper_001_receiver1_irq),            // interrupt_sender.irq
		.addr      (mm_interconnect_1_i2c_ext_csr_address),   //              csr.address
		.read      (mm_interconnect_1_i2c_ext_csr_read),      //                 .read
		.write     (mm_interconnect_1_i2c_ext_csr_write),     //                 .write
		.writedata (mm_interconnect_1_i2c_ext_csr_writedata), //                 .writedata
		.readdata  (mm_interconnect_1_i2c_ext_csr_readdata),  //                 .readdata
		.sda_in    (i2c_ext_sda_in),                          //       i2c_serial.sda_in
		.scl_in    (i2c_ext_scl_in),                          //                 .scl_in
		.sda_oe    (i2c_ext_sda_oe),                          //                 .sda_oe
		.scl_oe    (i2c_ext_scl_oe),                          //                 .scl_oe
		.src_data  (),                                        //      (terminated)
		.src_valid (),                                        //      (terminated)
		.src_ready (1'b0),                                    //      (terminated)
		.snk_data  (16'b0000000000000000),                    //      (terminated)
		.snk_valid (1'b0),                                    //      (terminated)
		.snk_ready ()                                         //      (terminated)
	);

	altera_avalon_i2c #(
		.USE_AV_ST       (0),
		.FIFO_DEPTH      (32),
		.FIFO_DEPTH_LOG2 (5)
	) i2c_int (
		.clk       (clk_clk),                                 //            clock.clk
		.rst_n     (~rst_controller_003_reset_out_reset),     //       reset_sink.reset_n
		.intr      (irq_mapper_001_receiver0_irq),            // interrupt_sender.irq
		.addr      (mm_interconnect_1_i2c_int_csr_address),   //              csr.address
		.read      (mm_interconnect_1_i2c_int_csr_read),      //                 .read
		.write     (mm_interconnect_1_i2c_int_csr_write),     //                 .write
		.writedata (mm_interconnect_1_i2c_int_csr_writedata), //                 .writedata
		.readdata  (mm_interconnect_1_i2c_int_csr_readdata),  //                 .readdata
		.sda_in    (i2c_int_sda_in),                          //       i2c_serial.sda_in
		.scl_in    (i2c_int_scl_in),                          //                 .scl_in
		.sda_oe    (i2c_int_sda_oe),                          //                 .sda_oe
		.scl_oe    (i2c_int_scl_oe),                          //                 .scl_oe
		.src_data  (),                                        //      (terminated)
		.src_valid (),                                        //      (terminated)
		.src_ready (1'b0),                                    //      (terminated)
		.snk_data  (16'b0000000000000000),                    //      (terminated)
		.snk_valid (1'b0),                                    //      (terminated)
		.snk_ready ()                                         //      (terminated)
	);

	soc_system_v5_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_003_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_1_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_1_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_1_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                   //               irq.irq
	);

	soc_system_v5_master_non_sec #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) master_non_sec (
		.clk_clk              (clk_clk),                             //          clk.clk
		.clk_reset_reset      (~reset_reset_n),                      //    clk_reset.reset
		.master_address       (master_non_sec_master_address),       //       master.address
		.master_readdata      (master_non_sec_master_readdata),      //             .readdata
		.master_read          (master_non_sec_master_read),          //             .read
		.master_write         (master_non_sec_master_write),         //             .write
		.master_writedata     (master_non_sec_master_writedata),     //             .writedata
		.master_waitrequest   (master_non_sec_master_waitrequest),   //             .waitrequest
		.master_readdatavalid (master_non_sec_master_readdatavalid), //             .readdatavalid
		.master_byteenable    (master_non_sec_master_byteenable),    //             .byteenable
		.master_reset_reset   ()                                     // master_reset.reset
	);

	soc_system_v5_master_non_sec #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) master_secure (
		.clk_clk              (clk_clk),                            //          clk.clk
		.clk_reset_reset      (~reset_reset_n),                     //    clk_reset.reset
		.master_address       (master_secure_master_address),       //       master.address
		.master_readdata      (master_secure_master_readdata),      //             .readdata
		.master_read          (master_secure_master_read),          //             .read
		.master_write         (master_secure_master_write),         //             .write
		.master_writedata     (master_secure_master_writedata),     //             .writedata
		.master_waitrequest   (master_secure_master_waitrequest),   //             .waitrequest
		.master_readdatavalid (master_secure_master_readdatavalid), //             .readdatavalid
		.master_byteenable    (master_secure_master_byteenable),    //             .byteenable
		.master_reset_reset   ()                                    // master_reset.reset
	);

	soc_system_v5_nmr_parameters nmr_parameters (
		.adc_val_sub_clk_clk                         (clk_clk),                                                         //                      adc_val_sub_clk.clk
		.adc_val_sub_external_connection_export      (adc_val_sub_export),                                              //      adc_val_sub_external_connection.export
		.adc_val_sub_reset_reset_n                   (~rst_controller_003_reset_out_reset),                             //                    adc_val_sub_reset.reset_n
		.adc_val_sub_s1_address                      (mm_interconnect_1_nmr_parameters_adc_val_sub_s1_address),         //                       adc_val_sub_s1.address
		.adc_val_sub_s1_write_n                      (~mm_interconnect_1_nmr_parameters_adc_val_sub_s1_write),          //                                     .write_n
		.adc_val_sub_s1_writedata                    (mm_interconnect_1_nmr_parameters_adc_val_sub_s1_writedata),       //                                     .writedata
		.adc_val_sub_s1_chipselect                   (mm_interconnect_1_nmr_parameters_adc_val_sub_s1_chipselect),      //                                     .chipselect
		.adc_val_sub_s1_readdata                     (mm_interconnect_1_nmr_parameters_adc_val_sub_s1_readdata),        //                                     .readdata
		.delay_nosig_clk_clk                         (clk_clk),                                                         //                      delay_nosig_clk.clk
		.delay_nosig_external_connection_export      (delay_nosig_export),                                              //      delay_nosig_external_connection.export
		.delay_nosig_reset_reset_n                   (~rst_controller_003_reset_out_reset),                             //                    delay_nosig_reset.reset_n
		.delay_nosig_s1_address                      (mm_interconnect_1_nmr_parameters_delay_nosig_s1_address),         //                       delay_nosig_s1.address
		.delay_nosig_s1_write_n                      (~mm_interconnect_1_nmr_parameters_delay_nosig_s1_write),          //                                     .write_n
		.delay_nosig_s1_writedata                    (mm_interconnect_1_nmr_parameters_delay_nosig_s1_writedata),       //                                     .writedata
		.delay_nosig_s1_chipselect                   (mm_interconnect_1_nmr_parameters_delay_nosig_s1_chipselect),      //                                     .chipselect
		.delay_nosig_s1_readdata                     (mm_interconnect_1_nmr_parameters_delay_nosig_s1_readdata),        //                                     .readdata
		.delay_sig_clk_clk                           (clk_clk),                                                         //                        delay_sig_clk.clk
		.delay_sig_external_connection_export        (delay_sig_export),                                                //        delay_sig_external_connection.export
		.delay_sig_reset_reset_n                     (~rst_controller_003_reset_out_reset),                             //                      delay_sig_reset.reset_n
		.delay_sig_s1_address                        (mm_interconnect_1_nmr_parameters_delay_sig_s1_address),           //                         delay_sig_s1.address
		.delay_sig_s1_write_n                        (~mm_interconnect_1_nmr_parameters_delay_sig_s1_write),            //                                     .write_n
		.delay_sig_s1_writedata                      (mm_interconnect_1_nmr_parameters_delay_sig_s1_writedata),         //                                     .writedata
		.delay_sig_s1_chipselect                     (mm_interconnect_1_nmr_parameters_delay_sig_s1_chipselect),        //                                     .chipselect
		.delay_sig_s1_readdata                       (mm_interconnect_1_nmr_parameters_delay_sig_s1_readdata),          //                                     .readdata
		.delay_t1_clk_clk                            (clk_clk),                                                         //                         delay_t1_clk.clk
		.delay_t1_external_connection_export         (delay_t1_export),                                                 //         delay_t1_external_connection.export
		.delay_t1_reset_reset_n                      (~rst_controller_003_reset_out_reset),                             //                       delay_t1_reset.reset_n
		.delay_t1_s1_address                         (mm_interconnect_1_nmr_parameters_delay_t1_s1_address),            //                          delay_t1_s1.address
		.delay_t1_s1_write_n                         (~mm_interconnect_1_nmr_parameters_delay_t1_s1_write),             //                                     .write_n
		.delay_t1_s1_writedata                       (mm_interconnect_1_nmr_parameters_delay_t1_s1_writedata),          //                                     .writedata
		.delay_t1_s1_chipselect                      (mm_interconnect_1_nmr_parameters_delay_t1_s1_chipselect),         //                                     .chipselect
		.delay_t1_s1_readdata                        (mm_interconnect_1_nmr_parameters_delay_t1_s1_readdata),           //                                     .readdata
		.echoes_per_scan_clk_clk                     (clk_clk),                                                         //                  echoes_per_scan_clk.clk
		.echoes_per_scan_external_connection_export  (echoes_per_scan_export),                                          //  echoes_per_scan_external_connection.export
		.echoes_per_scan_reset_reset_n               (~rst_controller_003_reset_out_reset),                             //                echoes_per_scan_reset.reset_n
		.echoes_per_scan_s1_address                  (mm_interconnect_1_nmr_parameters_echoes_per_scan_s1_address),     //                   echoes_per_scan_s1.address
		.echoes_per_scan_s1_write_n                  (~mm_interconnect_1_nmr_parameters_echoes_per_scan_s1_write),      //                                     .write_n
		.echoes_per_scan_s1_writedata                (mm_interconnect_1_nmr_parameters_echoes_per_scan_s1_writedata),   //                                     .writedata
		.echoes_per_scan_s1_chipselect               (mm_interconnect_1_nmr_parameters_echoes_per_scan_s1_chipselect),  //                                     .chipselect
		.echoes_per_scan_s1_readdata                 (mm_interconnect_1_nmr_parameters_echoes_per_scan_s1_readdata),    //                                     .readdata
		.init_delay_clk_clk                          (clk_clk),                                                         //                       init_delay_clk.clk
		.init_delay_external_connection_export       (init_delay_export),                                               //       init_delay_external_connection.export
		.init_delay_reset_reset_n                    (~rst_controller_003_reset_out_reset),                             //                     init_delay_reset.reset_n
		.init_delay_s1_address                       (mm_interconnect_1_nmr_parameters_init_delay_s1_address),          //                        init_delay_s1.address
		.init_delay_s1_write_n                       (~mm_interconnect_1_nmr_parameters_init_delay_s1_write),           //                                     .write_n
		.init_delay_s1_writedata                     (mm_interconnect_1_nmr_parameters_init_delay_s1_writedata),        //                                     .writedata
		.init_delay_s1_chipselect                    (mm_interconnect_1_nmr_parameters_init_delay_s1_chipselect),       //                                     .chipselect
		.init_delay_s1_readdata                      (mm_interconnect_1_nmr_parameters_init_delay_s1_readdata),         //                                     .readdata
		.pulse_180deg_clk_clk                        (clk_clk),                                                         //                     pulse_180deg_clk.clk
		.pulse_180deg_external_connection_export     (pulse_180deg_export),                                             //     pulse_180deg_external_connection.export
		.pulse_180deg_reset_reset_n                  (~rst_controller_003_reset_out_reset),                             //                   pulse_180deg_reset.reset_n
		.pulse_180deg_s1_address                     (mm_interconnect_1_nmr_parameters_pulse_180deg_s1_address),        //                      pulse_180deg_s1.address
		.pulse_180deg_s1_write_n                     (~mm_interconnect_1_nmr_parameters_pulse_180deg_s1_write),         //                                     .write_n
		.pulse_180deg_s1_writedata                   (mm_interconnect_1_nmr_parameters_pulse_180deg_s1_writedata),      //                                     .writedata
		.pulse_180deg_s1_chipselect                  (mm_interconnect_1_nmr_parameters_pulse_180deg_s1_chipselect),     //                                     .chipselect
		.pulse_180deg_s1_readdata                    (mm_interconnect_1_nmr_parameters_pulse_180deg_s1_readdata),       //                                     .readdata
		.pulse_90deg_clk_clk                         (clk_clk),                                                         //                      pulse_90deg_clk.clk
		.pulse_90deg_external_connection_export      (pulse_90deg_export),                                              //      pulse_90deg_external_connection.export
		.pulse_90deg_reset_reset_n                   (~rst_controller_003_reset_out_reset),                             //                    pulse_90deg_reset.reset_n
		.pulse_90deg_s1_address                      (mm_interconnect_1_nmr_parameters_pulse_90deg_s1_address),         //                       pulse_90deg_s1.address
		.pulse_90deg_s1_write_n                      (~mm_interconnect_1_nmr_parameters_pulse_90deg_s1_write),          //                                     .write_n
		.pulse_90deg_s1_writedata                    (mm_interconnect_1_nmr_parameters_pulse_90deg_s1_writedata),       //                                     .writedata
		.pulse_90deg_s1_chipselect                   (mm_interconnect_1_nmr_parameters_pulse_90deg_s1_chipselect),      //                                     .chipselect
		.pulse_90deg_s1_readdata                     (mm_interconnect_1_nmr_parameters_pulse_90deg_s1_readdata),        //                                     .readdata
		.pulse_t1_clk_clk                            (clk_clk),                                                         //                         pulse_t1_clk.clk
		.pulse_t1_external_connection_export         (pulse_t1_export),                                                 //         pulse_t1_external_connection.export
		.pulse_t1_reset_reset_n                      (~rst_controller_003_reset_out_reset),                             //                       pulse_t1_reset.reset_n
		.pulse_t1_s1_address                         (mm_interconnect_1_nmr_parameters_pulse_t1_s1_address),            //                          pulse_t1_s1.address
		.pulse_t1_s1_write_n                         (~mm_interconnect_1_nmr_parameters_pulse_t1_s1_write),             //                                     .write_n
		.pulse_t1_s1_writedata                       (mm_interconnect_1_nmr_parameters_pulse_t1_s1_writedata),          //                                     .writedata
		.pulse_t1_s1_chipselect                      (mm_interconnect_1_nmr_parameters_pulse_t1_s1_chipselect),         //                                     .chipselect
		.pulse_t1_s1_readdata                        (mm_interconnect_1_nmr_parameters_pulse_t1_s1_readdata),           //                                     .readdata
		.rx_delay_clk_clk                            (clk_clk),                                                         //                         rx_delay_clk.clk
		.rx_delay_external_connection_export         (rx_delay_export),                                                 //         rx_delay_external_connection.export
		.rx_delay_reset_reset_n                      (~rst_controller_003_reset_out_reset),                             //                       rx_delay_reset.reset_n
		.rx_delay_s1_address                         (mm_interconnect_1_nmr_parameters_rx_delay_s1_address),            //                          rx_delay_s1.address
		.rx_delay_s1_write_n                         (~mm_interconnect_1_nmr_parameters_rx_delay_s1_write),             //                                     .write_n
		.rx_delay_s1_writedata                       (mm_interconnect_1_nmr_parameters_rx_delay_s1_writedata),          //                                     .writedata
		.rx_delay_s1_chipselect                      (mm_interconnect_1_nmr_parameters_rx_delay_s1_chipselect),         //                                     .chipselect
		.rx_delay_s1_readdata                        (mm_interconnect_1_nmr_parameters_rx_delay_s1_readdata),           //                                     .readdata
		.samples_per_echo_clk_clk                    (clk_clk),                                                         //                 samples_per_echo_clk.clk
		.samples_per_echo_external_connection_export (samples_per_echo_export),                                         // samples_per_echo_external_connection.export
		.samples_per_echo_reset_reset_n              (~rst_controller_003_reset_out_reset),                             //               samples_per_echo_reset.reset_n
		.samples_per_echo_s1_address                 (mm_interconnect_1_nmr_parameters_samples_per_echo_s1_address),    //                  samples_per_echo_s1.address
		.samples_per_echo_s1_write_n                 (~mm_interconnect_1_nmr_parameters_samples_per_echo_s1_write),     //                                     .write_n
		.samples_per_echo_s1_writedata               (mm_interconnect_1_nmr_parameters_samples_per_echo_s1_writedata),  //                                     .writedata
		.samples_per_echo_s1_chipselect              (mm_interconnect_1_nmr_parameters_samples_per_echo_s1_chipselect), //                                     .chipselect
		.samples_per_echo_s1_readdata                (mm_interconnect_1_nmr_parameters_samples_per_echo_s1_readdata)    //                                     .readdata
	);

	soc_system_v5_nmr_sys_pll nmr_sys_pll (
		.refclk            (clk_clk),                                              //            refclk.clk
		.rst               (nmr_sys_pll_reset_reset),                              //             reset.reset
		.outclk_0          (nmr_sys_pll_outclk_clk),                               //           outclk0.clk
		.locked            (nmr_sys_pll_locked_export),                            //            locked.export
		.reconfig_to_pll   (nmr_sys_pll_reconfig_reconfig_to_pll_reconfig_to_pll), //   reconfig_to_pll.reconfig_to_pll
		.reconfig_from_pll (nmr_sys_pll_reconfig_from_pll_reconfig_from_pll)       // reconfig_from_pll.reconfig_from_pll
	);

	altera_pll_reconfig_top #(
		.device_family       ("Cyclone V"),
		.ENABLE_MIF          (0),
		.MIF_FILE_NAME       (""),
		.ENABLE_BYTEENABLE   (0),
		.BYTEENABLE_WIDTH    (4),
		.RECONFIG_ADDR_WIDTH (6),
		.RECONFIG_DATA_WIDTH (32),
		.reconf_width        (64),
		.WAIT_FOR_LOCK       (1)
	) nmr_sys_pll_reconfig (
		.mgmt_clk          (clk_clk),                                                              //          mgmt_clk.clk
		.mgmt_reset        (rst_controller_003_reset_out_reset),                                   //        mgmt_reset.reset
		.mgmt_waitrequest  (mm_interconnect_1_nmr_sys_pll_reconfig_mgmt_avalon_slave_waitrequest), // mgmt_avalon_slave.waitrequest
		.mgmt_read         (mm_interconnect_1_nmr_sys_pll_reconfig_mgmt_avalon_slave_read),        //                  .read
		.mgmt_write        (mm_interconnect_1_nmr_sys_pll_reconfig_mgmt_avalon_slave_write),       //                  .write
		.mgmt_readdata     (mm_interconnect_1_nmr_sys_pll_reconfig_mgmt_avalon_slave_readdata),    //                  .readdata
		.mgmt_address      (mm_interconnect_1_nmr_sys_pll_reconfig_mgmt_avalon_slave_address),     //                  .address
		.mgmt_writedata    (mm_interconnect_1_nmr_sys_pll_reconfig_mgmt_avalon_slave_writedata),   //                  .writedata
		.reconfig_to_pll   (nmr_sys_pll_reconfig_reconfig_to_pll_reconfig_to_pll),                 //   reconfig_to_pll.reconfig_to_pll
		.reconfig_from_pll (nmr_sys_pll_reconfig_from_pll_reconfig_from_pll),                      // reconfig_from_pll.reconfig_from_pll
		.mgmt_byteenable   (4'b0000)                                                               //       (terminated)
	);

	soc_system_v5_sdram sdram (
		.clk            (clk_clk),                                  //   clk.clk
		.reset_n        (~rst_controller_003_reset_out_reset),      // reset.reset_n
		.az_addr        (mm_interconnect_1_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_1_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_1_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_1_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_1_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_1_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_1_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_1_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_1_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	soc_system_v5_spi_afe_relays spi_afe_relays (
		.clk           (clk_clk),                                                      //              clk.clk
		.reset_n       (~rst_controller_003_reset_out_reset),                          //            reset.reset_n
		.data_from_cpu (mm_interconnect_1_spi_afe_relays_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_1_spi_afe_relays_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_1_spi_afe_relays_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_1_spi_afe_relays_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_1_spi_afe_relays_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_1_spi_afe_relays_spi_control_port_write),     //                 .write_n
		.irq           (irq_mapper_001_receiver7_irq),                                 //              irq.irq
		.MISO          (spi_afe_relays_MISO),                                          //         external.export
		.MOSI          (spi_afe_relays_MOSI),                                          //                 .export
		.SCLK          (spi_afe_relays_SCLK),                                          //                 .export
		.SS_n          (spi_afe_relays_SS_n)                                           //                 .export
	);

	soc_system_v5_spi_afe_relays spi_mtch_ntwrk (
		.clk           (clk_clk),                                                      //              clk.clk
		.reset_n       (~rst_controller_003_reset_out_reset),                          //            reset.reset_n
		.data_from_cpu (mm_interconnect_1_spi_mtch_ntwrk_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_1_spi_mtch_ntwrk_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_1_spi_mtch_ntwrk_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_1_spi_mtch_ntwrk_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_1_spi_mtch_ntwrk_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_1_spi_mtch_ntwrk_spi_control_port_write),     //                 .write_n
		.irq           (irq_mapper_001_receiver4_irq),                                 //              irq.irq
		.MISO          (spi_mtch_ntwrk_MISO),                                          //         external.export
		.MOSI          (spi_mtch_ntwrk_MOSI),                                          //                 .export
		.SCLK          (spi_mtch_ntwrk_SCLK),                                          //                 .export
		.SS_n          (spi_mtch_ntwrk_SS_n)                                           //                 .export
	);

	soc_system_v5_switches switches (
		.clk      (clk_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_003_reset_out_reset),    //               reset.reset_n
		.address  (mm_interconnect_1_switches_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_switches_s1_readdata), //                    .readdata
		.in_port  (switches_export)                         // external_connection.export
	);

	soc_system_v5_sysid_qsys sysid_qsys (
		.clock    (clk_clk),                                             //           clk.clk
		.reset_n  (~rst_controller_003_reset_out_reset),                 //         reset.reset_n
		.readdata (mm_interconnect_1_sysid_qsys_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_1_sysid_qsys_control_slave_address)   //              .address
	);

	soc_system_v5_mm_interconnect_0 mm_interconnect_0 (
		.hps_0_f2h_axi_slave_awid                                         (mm_interconnect_0_hps_0_f2h_axi_slave_awid),    //                                        hps_0_f2h_axi_slave.awid
		.hps_0_f2h_axi_slave_awaddr                                       (mm_interconnect_0_hps_0_f2h_axi_slave_awaddr),  //                                                           .awaddr
		.hps_0_f2h_axi_slave_awlen                                        (mm_interconnect_0_hps_0_f2h_axi_slave_awlen),   //                                                           .awlen
		.hps_0_f2h_axi_slave_awsize                                       (mm_interconnect_0_hps_0_f2h_axi_slave_awsize),  //                                                           .awsize
		.hps_0_f2h_axi_slave_awburst                                      (mm_interconnect_0_hps_0_f2h_axi_slave_awburst), //                                                           .awburst
		.hps_0_f2h_axi_slave_awlock                                       (mm_interconnect_0_hps_0_f2h_axi_slave_awlock),  //                                                           .awlock
		.hps_0_f2h_axi_slave_awcache                                      (mm_interconnect_0_hps_0_f2h_axi_slave_awcache), //                                                           .awcache
		.hps_0_f2h_axi_slave_awprot                                       (mm_interconnect_0_hps_0_f2h_axi_slave_awprot),  //                                                           .awprot
		.hps_0_f2h_axi_slave_awuser                                       (mm_interconnect_0_hps_0_f2h_axi_slave_awuser),  //                                                           .awuser
		.hps_0_f2h_axi_slave_awvalid                                      (mm_interconnect_0_hps_0_f2h_axi_slave_awvalid), //                                                           .awvalid
		.hps_0_f2h_axi_slave_awready                                      (mm_interconnect_0_hps_0_f2h_axi_slave_awready), //                                                           .awready
		.hps_0_f2h_axi_slave_wid                                          (mm_interconnect_0_hps_0_f2h_axi_slave_wid),     //                                                           .wid
		.hps_0_f2h_axi_slave_wdata                                        (mm_interconnect_0_hps_0_f2h_axi_slave_wdata),   //                                                           .wdata
		.hps_0_f2h_axi_slave_wstrb                                        (mm_interconnect_0_hps_0_f2h_axi_slave_wstrb),   //                                                           .wstrb
		.hps_0_f2h_axi_slave_wlast                                        (mm_interconnect_0_hps_0_f2h_axi_slave_wlast),   //                                                           .wlast
		.hps_0_f2h_axi_slave_wvalid                                       (mm_interconnect_0_hps_0_f2h_axi_slave_wvalid),  //                                                           .wvalid
		.hps_0_f2h_axi_slave_wready                                       (mm_interconnect_0_hps_0_f2h_axi_slave_wready),  //                                                           .wready
		.hps_0_f2h_axi_slave_bid                                          (mm_interconnect_0_hps_0_f2h_axi_slave_bid),     //                                                           .bid
		.hps_0_f2h_axi_slave_bresp                                        (mm_interconnect_0_hps_0_f2h_axi_slave_bresp),   //                                                           .bresp
		.hps_0_f2h_axi_slave_bvalid                                       (mm_interconnect_0_hps_0_f2h_axi_slave_bvalid),  //                                                           .bvalid
		.hps_0_f2h_axi_slave_bready                                       (mm_interconnect_0_hps_0_f2h_axi_slave_bready),  //                                                           .bready
		.hps_0_f2h_axi_slave_arid                                         (mm_interconnect_0_hps_0_f2h_axi_slave_arid),    //                                                           .arid
		.hps_0_f2h_axi_slave_araddr                                       (mm_interconnect_0_hps_0_f2h_axi_slave_araddr),  //                                                           .araddr
		.hps_0_f2h_axi_slave_arlen                                        (mm_interconnect_0_hps_0_f2h_axi_slave_arlen),   //                                                           .arlen
		.hps_0_f2h_axi_slave_arsize                                       (mm_interconnect_0_hps_0_f2h_axi_slave_arsize),  //                                                           .arsize
		.hps_0_f2h_axi_slave_arburst                                      (mm_interconnect_0_hps_0_f2h_axi_slave_arburst), //                                                           .arburst
		.hps_0_f2h_axi_slave_arlock                                       (mm_interconnect_0_hps_0_f2h_axi_slave_arlock),  //                                                           .arlock
		.hps_0_f2h_axi_slave_arcache                                      (mm_interconnect_0_hps_0_f2h_axi_slave_arcache), //                                                           .arcache
		.hps_0_f2h_axi_slave_arprot                                       (mm_interconnect_0_hps_0_f2h_axi_slave_arprot),  //                                                           .arprot
		.hps_0_f2h_axi_slave_aruser                                       (mm_interconnect_0_hps_0_f2h_axi_slave_aruser),  //                                                           .aruser
		.hps_0_f2h_axi_slave_arvalid                                      (mm_interconnect_0_hps_0_f2h_axi_slave_arvalid), //                                                           .arvalid
		.hps_0_f2h_axi_slave_arready                                      (mm_interconnect_0_hps_0_f2h_axi_slave_arready), //                                                           .arready
		.hps_0_f2h_axi_slave_rid                                          (mm_interconnect_0_hps_0_f2h_axi_slave_rid),     //                                                           .rid
		.hps_0_f2h_axi_slave_rdata                                        (mm_interconnect_0_hps_0_f2h_axi_slave_rdata),   //                                                           .rdata
		.hps_0_f2h_axi_slave_rresp                                        (mm_interconnect_0_hps_0_f2h_axi_slave_rresp),   //                                                           .rresp
		.hps_0_f2h_axi_slave_rlast                                        (mm_interconnect_0_hps_0_f2h_axi_slave_rlast),   //                                                           .rlast
		.hps_0_f2h_axi_slave_rvalid                                       (mm_interconnect_0_hps_0_f2h_axi_slave_rvalid),  //                                                           .rvalid
		.hps_0_f2h_axi_slave_rready                                       (mm_interconnect_0_hps_0_f2h_axi_slave_rready),  //                                                           .rready
		.clk_0_clk_clk                                                    (clk_clk),                                       //                                                  clk_0_clk.clk
		.alt_vip_vfr_vga_clock_master_reset_reset_bridge_in_reset_reset   (rst_controller_003_reset_out_reset),            //   alt_vip_vfr_vga_clock_master_reset_reset_bridge_in_reset.reset
		.hps_0_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset_reset (rst_controller_004_reset_out_reset),            // hps_0_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset.reset
		.master_secure_clk_reset_reset_bridge_in_reset_reset              (rst_controller_003_reset_out_reset),            //              master_secure_clk_reset_reset_bridge_in_reset.reset
		.alt_vip_vfr_vga_avalon_master_address                            (alt_vip_vfr_vga_avalon_master_address),         //                              alt_vip_vfr_vga_avalon_master.address
		.alt_vip_vfr_vga_avalon_master_waitrequest                        (alt_vip_vfr_vga_avalon_master_waitrequest),     //                                                           .waitrequest
		.alt_vip_vfr_vga_avalon_master_burstcount                         (alt_vip_vfr_vga_avalon_master_burstcount),      //                                                           .burstcount
		.alt_vip_vfr_vga_avalon_master_read                               (alt_vip_vfr_vga_avalon_master_read),            //                                                           .read
		.alt_vip_vfr_vga_avalon_master_readdata                           (alt_vip_vfr_vga_avalon_master_readdata),        //                                                           .readdata
		.alt_vip_vfr_vga_avalon_master_readdatavalid                      (alt_vip_vfr_vga_avalon_master_readdatavalid),   //                                                           .readdatavalid
		.master_secure_master_address                                     (master_secure_master_address),                  //                                       master_secure_master.address
		.master_secure_master_waitrequest                                 (master_secure_master_waitrequest),              //                                                           .waitrequest
		.master_secure_master_byteenable                                  (master_secure_master_byteenable),               //                                                           .byteenable
		.master_secure_master_read                                        (master_secure_master_read),                     //                                                           .read
		.master_secure_master_readdata                                    (master_secure_master_readdata),                 //                                                           .readdata
		.master_secure_master_readdatavalid                               (master_secure_master_readdatavalid),            //                                                           .readdatavalid
		.master_secure_master_write                                       (master_secure_master_write),                    //                                                           .write
		.master_secure_master_writedata                                   (master_secure_master_writedata)                 //                                                           .writedata
	);

	soc_system_v5_mm_interconnect_1 mm_interconnect_1 (
		.hps_0_h2f_axi_master_awid                                        (hps_0_h2f_axi_master_awid),                                             //                                       hps_0_h2f_axi_master.awid
		.hps_0_h2f_axi_master_awaddr                                      (hps_0_h2f_axi_master_awaddr),                                           //                                                           .awaddr
		.hps_0_h2f_axi_master_awlen                                       (hps_0_h2f_axi_master_awlen),                                            //                                                           .awlen
		.hps_0_h2f_axi_master_awsize                                      (hps_0_h2f_axi_master_awsize),                                           //                                                           .awsize
		.hps_0_h2f_axi_master_awburst                                     (hps_0_h2f_axi_master_awburst),                                          //                                                           .awburst
		.hps_0_h2f_axi_master_awlock                                      (hps_0_h2f_axi_master_awlock),                                           //                                                           .awlock
		.hps_0_h2f_axi_master_awcache                                     (hps_0_h2f_axi_master_awcache),                                          //                                                           .awcache
		.hps_0_h2f_axi_master_awprot                                      (hps_0_h2f_axi_master_awprot),                                           //                                                           .awprot
		.hps_0_h2f_axi_master_awvalid                                     (hps_0_h2f_axi_master_awvalid),                                          //                                                           .awvalid
		.hps_0_h2f_axi_master_awready                                     (hps_0_h2f_axi_master_awready),                                          //                                                           .awready
		.hps_0_h2f_axi_master_wid                                         (hps_0_h2f_axi_master_wid),                                              //                                                           .wid
		.hps_0_h2f_axi_master_wdata                                       (hps_0_h2f_axi_master_wdata),                                            //                                                           .wdata
		.hps_0_h2f_axi_master_wstrb                                       (hps_0_h2f_axi_master_wstrb),                                            //                                                           .wstrb
		.hps_0_h2f_axi_master_wlast                                       (hps_0_h2f_axi_master_wlast),                                            //                                                           .wlast
		.hps_0_h2f_axi_master_wvalid                                      (hps_0_h2f_axi_master_wvalid),                                           //                                                           .wvalid
		.hps_0_h2f_axi_master_wready                                      (hps_0_h2f_axi_master_wready),                                           //                                                           .wready
		.hps_0_h2f_axi_master_bid                                         (hps_0_h2f_axi_master_bid),                                              //                                                           .bid
		.hps_0_h2f_axi_master_bresp                                       (hps_0_h2f_axi_master_bresp),                                            //                                                           .bresp
		.hps_0_h2f_axi_master_bvalid                                      (hps_0_h2f_axi_master_bvalid),                                           //                                                           .bvalid
		.hps_0_h2f_axi_master_bready                                      (hps_0_h2f_axi_master_bready),                                           //                                                           .bready
		.hps_0_h2f_axi_master_arid                                        (hps_0_h2f_axi_master_arid),                                             //                                                           .arid
		.hps_0_h2f_axi_master_araddr                                      (hps_0_h2f_axi_master_araddr),                                           //                                                           .araddr
		.hps_0_h2f_axi_master_arlen                                       (hps_0_h2f_axi_master_arlen),                                            //                                                           .arlen
		.hps_0_h2f_axi_master_arsize                                      (hps_0_h2f_axi_master_arsize),                                           //                                                           .arsize
		.hps_0_h2f_axi_master_arburst                                     (hps_0_h2f_axi_master_arburst),                                          //                                                           .arburst
		.hps_0_h2f_axi_master_arlock                                      (hps_0_h2f_axi_master_arlock),                                           //                                                           .arlock
		.hps_0_h2f_axi_master_arcache                                     (hps_0_h2f_axi_master_arcache),                                          //                                                           .arcache
		.hps_0_h2f_axi_master_arprot                                      (hps_0_h2f_axi_master_arprot),                                           //                                                           .arprot
		.hps_0_h2f_axi_master_arvalid                                     (hps_0_h2f_axi_master_arvalid),                                          //                                                           .arvalid
		.hps_0_h2f_axi_master_arready                                     (hps_0_h2f_axi_master_arready),                                          //                                                           .arready
		.hps_0_h2f_axi_master_rid                                         (hps_0_h2f_axi_master_rid),                                              //                                                           .rid
		.hps_0_h2f_axi_master_rdata                                       (hps_0_h2f_axi_master_rdata),                                            //                                                           .rdata
		.hps_0_h2f_axi_master_rresp                                       (hps_0_h2f_axi_master_rresp),                                            //                                                           .rresp
		.hps_0_h2f_axi_master_rlast                                       (hps_0_h2f_axi_master_rlast),                                            //                                                           .rlast
		.hps_0_h2f_axi_master_rvalid                                      (hps_0_h2f_axi_master_rvalid),                                           //                                                           .rvalid
		.hps_0_h2f_axi_master_rready                                      (hps_0_h2f_axi_master_rready),                                           //                                                           .rready
		.hps_0_h2f_lw_axi_master_awid                                     (hps_0_h2f_lw_axi_master_awid),                                          //                                    hps_0_h2f_lw_axi_master.awid
		.hps_0_h2f_lw_axi_master_awaddr                                   (hps_0_h2f_lw_axi_master_awaddr),                                        //                                                           .awaddr
		.hps_0_h2f_lw_axi_master_awlen                                    (hps_0_h2f_lw_axi_master_awlen),                                         //                                                           .awlen
		.hps_0_h2f_lw_axi_master_awsize                                   (hps_0_h2f_lw_axi_master_awsize),                                        //                                                           .awsize
		.hps_0_h2f_lw_axi_master_awburst                                  (hps_0_h2f_lw_axi_master_awburst),                                       //                                                           .awburst
		.hps_0_h2f_lw_axi_master_awlock                                   (hps_0_h2f_lw_axi_master_awlock),                                        //                                                           .awlock
		.hps_0_h2f_lw_axi_master_awcache                                  (hps_0_h2f_lw_axi_master_awcache),                                       //                                                           .awcache
		.hps_0_h2f_lw_axi_master_awprot                                   (hps_0_h2f_lw_axi_master_awprot),                                        //                                                           .awprot
		.hps_0_h2f_lw_axi_master_awvalid                                  (hps_0_h2f_lw_axi_master_awvalid),                                       //                                                           .awvalid
		.hps_0_h2f_lw_axi_master_awready                                  (hps_0_h2f_lw_axi_master_awready),                                       //                                                           .awready
		.hps_0_h2f_lw_axi_master_wid                                      (hps_0_h2f_lw_axi_master_wid),                                           //                                                           .wid
		.hps_0_h2f_lw_axi_master_wdata                                    (hps_0_h2f_lw_axi_master_wdata),                                         //                                                           .wdata
		.hps_0_h2f_lw_axi_master_wstrb                                    (hps_0_h2f_lw_axi_master_wstrb),                                         //                                                           .wstrb
		.hps_0_h2f_lw_axi_master_wlast                                    (hps_0_h2f_lw_axi_master_wlast),                                         //                                                           .wlast
		.hps_0_h2f_lw_axi_master_wvalid                                   (hps_0_h2f_lw_axi_master_wvalid),                                        //                                                           .wvalid
		.hps_0_h2f_lw_axi_master_wready                                   (hps_0_h2f_lw_axi_master_wready),                                        //                                                           .wready
		.hps_0_h2f_lw_axi_master_bid                                      (hps_0_h2f_lw_axi_master_bid),                                           //                                                           .bid
		.hps_0_h2f_lw_axi_master_bresp                                    (hps_0_h2f_lw_axi_master_bresp),                                         //                                                           .bresp
		.hps_0_h2f_lw_axi_master_bvalid                                   (hps_0_h2f_lw_axi_master_bvalid),                                        //                                                           .bvalid
		.hps_0_h2f_lw_axi_master_bready                                   (hps_0_h2f_lw_axi_master_bready),                                        //                                                           .bready
		.hps_0_h2f_lw_axi_master_arid                                     (hps_0_h2f_lw_axi_master_arid),                                          //                                                           .arid
		.hps_0_h2f_lw_axi_master_araddr                                   (hps_0_h2f_lw_axi_master_araddr),                                        //                                                           .araddr
		.hps_0_h2f_lw_axi_master_arlen                                    (hps_0_h2f_lw_axi_master_arlen),                                         //                                                           .arlen
		.hps_0_h2f_lw_axi_master_arsize                                   (hps_0_h2f_lw_axi_master_arsize),                                        //                                                           .arsize
		.hps_0_h2f_lw_axi_master_arburst                                  (hps_0_h2f_lw_axi_master_arburst),                                       //                                                           .arburst
		.hps_0_h2f_lw_axi_master_arlock                                   (hps_0_h2f_lw_axi_master_arlock),                                        //                                                           .arlock
		.hps_0_h2f_lw_axi_master_arcache                                  (hps_0_h2f_lw_axi_master_arcache),                                       //                                                           .arcache
		.hps_0_h2f_lw_axi_master_arprot                                   (hps_0_h2f_lw_axi_master_arprot),                                        //                                                           .arprot
		.hps_0_h2f_lw_axi_master_arvalid                                  (hps_0_h2f_lw_axi_master_arvalid),                                       //                                                           .arvalid
		.hps_0_h2f_lw_axi_master_arready                                  (hps_0_h2f_lw_axi_master_arready),                                       //                                                           .arready
		.hps_0_h2f_lw_axi_master_rid                                      (hps_0_h2f_lw_axi_master_rid),                                           //                                                           .rid
		.hps_0_h2f_lw_axi_master_rdata                                    (hps_0_h2f_lw_axi_master_rdata),                                         //                                                           .rdata
		.hps_0_h2f_lw_axi_master_rresp                                    (hps_0_h2f_lw_axi_master_rresp),                                         //                                                           .rresp
		.hps_0_h2f_lw_axi_master_rlast                                    (hps_0_h2f_lw_axi_master_rlast),                                         //                                                           .rlast
		.hps_0_h2f_lw_axi_master_rvalid                                   (hps_0_h2f_lw_axi_master_rvalid),                                        //                                                           .rvalid
		.hps_0_h2f_lw_axi_master_rready                                   (hps_0_h2f_lw_axi_master_rready),                                        //                                                           .rready
		.clk_0_clk_clk                                                    (clk_clk),                                                               //                                                  clk_0_clk.clk
		.gp_pll_outclk0_clk                                               (gp_pll_outclk0_clk),                                                    //                                             gp_pll_outclk0.clk
		.adc_fifo_mem_reset_in_reset_bridge_in_reset_reset                (rst_controller_001_reset_out_reset),                                    //                adc_fifo_mem_reset_in_reset_bridge_in_reset.reset
		.alt_vip_vfr_vga_clock_reset_reset_reset_bridge_in_reset_reset    (rst_controller_002_reset_out_reset),                                    //    alt_vip_vfr_vga_clock_reset_reset_reset_bridge_in_reset.reset
		.dma_fifo_reset_reset_bridge_in_reset_reset                       (rst_controller_003_reset_out_reset),                                    //                       dma_fifo_reset_reset_bridge_in_reset.reset
		.hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_004_reset_out_reset),                                    // hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.master_non_sec_clk_reset_reset_bridge_in_reset_reset             (rst_controller_003_reset_out_reset),                                    //             master_non_sec_clk_reset_reset_bridge_in_reset.reset
		.dma_dconvi_read_master_address                                   (dma_dconvi_read_master_address),                                        //                                     dma_dconvi_read_master.address
		.dma_dconvi_read_master_waitrequest                               (dma_dconvi_read_master_waitrequest),                                    //                                                           .waitrequest
		.dma_dconvi_read_master_chipselect                                (dma_dconvi_read_master_chipselect),                                     //                                                           .chipselect
		.dma_dconvi_read_master_read                                      (~dma_dconvi_read_master_read),                                          //                                                           .read
		.dma_dconvi_read_master_readdata                                  (dma_dconvi_read_master_readdata),                                       //                                                           .readdata
		.dma_dconvi_read_master_readdatavalid                             (dma_dconvi_read_master_readdatavalid),                                  //                                                           .readdatavalid
		.dma_dconvi_write_master_address                                  (dma_dconvi_write_master_address),                                       //                                    dma_dconvi_write_master.address
		.dma_dconvi_write_master_waitrequest                              (dma_dconvi_write_master_waitrequest),                                   //                                                           .waitrequest
		.dma_dconvi_write_master_byteenable                               (dma_dconvi_write_master_byteenable),                                    //                                                           .byteenable
		.dma_dconvi_write_master_chipselect                               (dma_dconvi_write_master_chipselect),                                    //                                                           .chipselect
		.dma_dconvi_write_master_write                                    (~dma_dconvi_write_master_write),                                        //                                                           .write
		.dma_dconvi_write_master_writedata                                (dma_dconvi_write_master_writedata),                                     //                                                           .writedata
		.dma_dconvq_read_master_address                                   (dma_dconvq_read_master_address),                                        //                                     dma_dconvq_read_master.address
		.dma_dconvq_read_master_waitrequest                               (dma_dconvq_read_master_waitrequest),                                    //                                                           .waitrequest
		.dma_dconvq_read_master_chipselect                                (dma_dconvq_read_master_chipselect),                                     //                                                           .chipselect
		.dma_dconvq_read_master_read                                      (~dma_dconvq_read_master_read),                                          //                                                           .read
		.dma_dconvq_read_master_readdata                                  (dma_dconvq_read_master_readdata),                                       //                                                           .readdata
		.dma_dconvq_read_master_readdatavalid                             (dma_dconvq_read_master_readdatavalid),                                  //                                                           .readdatavalid
		.dma_dconvq_write_master_address                                  (dma_dconvq_write_master_address),                                       //                                    dma_dconvq_write_master.address
		.dma_dconvq_write_master_waitrequest                              (dma_dconvq_write_master_waitrequest),                                   //                                                           .waitrequest
		.dma_dconvq_write_master_byteenable                               (dma_dconvq_write_master_byteenable),                                    //                                                           .byteenable
		.dma_dconvq_write_master_chipselect                               (dma_dconvq_write_master_chipselect),                                    //                                                           .chipselect
		.dma_dconvq_write_master_write                                    (~dma_dconvq_write_master_write),                                        //                                                           .write
		.dma_dconvq_write_master_writedata                                (dma_dconvq_write_master_writedata),                                     //                                                           .writedata
		.dma_dummy_read_master_address                                    (dma_dummy_read_master_address),                                         //                                      dma_dummy_read_master.address
		.dma_dummy_read_master_waitrequest                                (dma_dummy_read_master_waitrequest),                                     //                                                           .waitrequest
		.dma_dummy_read_master_chipselect                                 (dma_dummy_read_master_chipselect),                                      //                                                           .chipselect
		.dma_dummy_read_master_read                                       (~dma_dummy_read_master_read),                                           //                                                           .read
		.dma_dummy_read_master_readdata                                   (dma_dummy_read_master_readdata),                                        //                                                           .readdata
		.dma_dummy_read_master_readdatavalid                              (dma_dummy_read_master_readdatavalid),                                   //                                                           .readdatavalid
		.dma_dummy_write_master_address                                   (dma_dummy_write_master_address),                                        //                                     dma_dummy_write_master.address
		.dma_dummy_write_master_waitrequest                               (dma_dummy_write_master_waitrequest),                                    //                                                           .waitrequest
		.dma_dummy_write_master_byteenable                                (dma_dummy_write_master_byteenable),                                     //                                                           .byteenable
		.dma_dummy_write_master_chipselect                                (dma_dummy_write_master_chipselect),                                     //                                                           .chipselect
		.dma_dummy_write_master_write                                     (~dma_dummy_write_master_write),                                         //                                                           .write
		.dma_dummy_write_master_writedata                                 (dma_dummy_write_master_writedata),                                      //                                                           .writedata
		.dma_fifo_read_master_address                                     (dma_fifo_read_master_address),                                          //                                       dma_fifo_read_master.address
		.dma_fifo_read_master_waitrequest                                 (dma_fifo_read_master_waitrequest),                                      //                                                           .waitrequest
		.dma_fifo_read_master_chipselect                                  (dma_fifo_read_master_chipselect),                                       //                                                           .chipselect
		.dma_fifo_read_master_read                                        (~dma_fifo_read_master_read),                                            //                                                           .read
		.dma_fifo_read_master_readdata                                    (dma_fifo_read_master_readdata),                                         //                                                           .readdata
		.dma_fifo_read_master_readdatavalid                               (dma_fifo_read_master_readdatavalid),                                    //                                                           .readdatavalid
		.dma_fifo_write_master_address                                    (dma_fifo_write_master_address),                                         //                                      dma_fifo_write_master.address
		.dma_fifo_write_master_waitrequest                                (dma_fifo_write_master_waitrequest),                                     //                                                           .waitrequest
		.dma_fifo_write_master_byteenable                                 (dma_fifo_write_master_byteenable),                                      //                                                           .byteenable
		.dma_fifo_write_master_chipselect                                 (dma_fifo_write_master_chipselect),                                      //                                                           .chipselect
		.dma_fifo_write_master_write                                      (~dma_fifo_write_master_write),                                          //                                                           .write
		.dma_fifo_write_master_writedata                                  (dma_fifo_write_master_writedata),                                       //                                                           .writedata
		.master_non_sec_master_address                                    (master_non_sec_master_address),                                         //                                      master_non_sec_master.address
		.master_non_sec_master_waitrequest                                (master_non_sec_master_waitrequest),                                     //                                                           .waitrequest
		.master_non_sec_master_byteenable                                 (master_non_sec_master_byteenable),                                      //                                                           .byteenable
		.master_non_sec_master_read                                       (master_non_sec_master_read),                                            //                                                           .read
		.master_non_sec_master_readdata                                   (master_non_sec_master_readdata),                                        //                                                           .readdata
		.master_non_sec_master_readdatavalid                              (master_non_sec_master_readdatavalid),                                   //                                                           .readdatavalid
		.master_non_sec_master_write                                      (master_non_sec_master_write),                                           //                                                           .write
		.master_non_sec_master_writedata                                  (master_non_sec_master_writedata),                                       //                                                           .writedata
		.adc_fifo_mem_in_csr_address                                      (mm_interconnect_1_adc_fifo_mem_in_csr_address),                         //                                        adc_fifo_mem_in_csr.address
		.adc_fifo_mem_in_csr_write                                        (mm_interconnect_1_adc_fifo_mem_in_csr_write),                           //                                                           .write
		.adc_fifo_mem_in_csr_read                                         (mm_interconnect_1_adc_fifo_mem_in_csr_read),                            //                                                           .read
		.adc_fifo_mem_in_csr_readdata                                     (mm_interconnect_1_adc_fifo_mem_in_csr_readdata),                        //                                                           .readdata
		.adc_fifo_mem_in_csr_writedata                                    (mm_interconnect_1_adc_fifo_mem_in_csr_writedata),                       //                                                           .writedata
		.adc_fifo_mem_out_address                                         (mm_interconnect_1_adc_fifo_mem_out_address),                            //                                           adc_fifo_mem_out.address
		.adc_fifo_mem_out_read                                            (mm_interconnect_1_adc_fifo_mem_out_read),                               //                                                           .read
		.adc_fifo_mem_out_readdata                                        (mm_interconnect_1_adc_fifo_mem_out_readdata),                           //                                                           .readdata
		.adc_fifo_mem_out_waitrequest                                     (mm_interconnect_1_adc_fifo_mem_out_waitrequest),                        //                                                           .waitrequest
		.alt_vip_vfr_vga_avalon_slave_address                             (mm_interconnect_1_alt_vip_vfr_vga_avalon_slave_address),                //                               alt_vip_vfr_vga_avalon_slave.address
		.alt_vip_vfr_vga_avalon_slave_write                               (mm_interconnect_1_alt_vip_vfr_vga_avalon_slave_write),                  //                                                           .write
		.alt_vip_vfr_vga_avalon_slave_read                                (mm_interconnect_1_alt_vip_vfr_vga_avalon_slave_read),                   //                                                           .read
		.alt_vip_vfr_vga_avalon_slave_readdata                            (mm_interconnect_1_alt_vip_vfr_vga_avalon_slave_readdata),               //                                                           .readdata
		.alt_vip_vfr_vga_avalon_slave_writedata                           (mm_interconnect_1_alt_vip_vfr_vga_avalon_slave_writedata),              //                                                           .writedata
		.analyzer_pll_reconfig_mgmt_avalon_slave_address                  (mm_interconnect_1_analyzer_pll_reconfig_mgmt_avalon_slave_address),     //                    analyzer_pll_reconfig_mgmt_avalon_slave.address
		.analyzer_pll_reconfig_mgmt_avalon_slave_write                    (mm_interconnect_1_analyzer_pll_reconfig_mgmt_avalon_slave_write),       //                                                           .write
		.analyzer_pll_reconfig_mgmt_avalon_slave_read                     (mm_interconnect_1_analyzer_pll_reconfig_mgmt_avalon_slave_read),        //                                                           .read
		.analyzer_pll_reconfig_mgmt_avalon_slave_readdata                 (mm_interconnect_1_analyzer_pll_reconfig_mgmt_avalon_slave_readdata),    //                                                           .readdata
		.analyzer_pll_reconfig_mgmt_avalon_slave_writedata                (mm_interconnect_1_analyzer_pll_reconfig_mgmt_avalon_slave_writedata),   //                                                           .writedata
		.analyzer_pll_reconfig_mgmt_avalon_slave_waitrequest              (mm_interconnect_1_analyzer_pll_reconfig_mgmt_avalon_slave_waitrequest), //                                                           .waitrequest
		.aux_cnt_out_s1_address                                           (mm_interconnect_1_aux_cnt_out_s1_address),                              //                                             aux_cnt_out_s1.address
		.aux_cnt_out_s1_write                                             (mm_interconnect_1_aux_cnt_out_s1_write),                                //                                                           .write
		.aux_cnt_out_s1_readdata                                          (mm_interconnect_1_aux_cnt_out_s1_readdata),                             //                                                           .readdata
		.aux_cnt_out_s1_writedata                                         (mm_interconnect_1_aux_cnt_out_s1_writedata),                            //                                                           .writedata
		.aux_cnt_out_s1_chipselect                                        (mm_interconnect_1_aux_cnt_out_s1_chipselect),                           //                                                           .chipselect
		.ctrl_in_s1_address                                               (mm_interconnect_1_ctrl_in_s1_address),                                  //                                                 ctrl_in_s1.address
		.ctrl_in_s1_readdata                                              (mm_interconnect_1_ctrl_in_s1_readdata),                                 //                                                           .readdata
		.ctrl_out_s1_address                                              (mm_interconnect_1_ctrl_out_s1_address),                                 //                                                ctrl_out_s1.address
		.ctrl_out_s1_write                                                (mm_interconnect_1_ctrl_out_s1_write),                                   //                                                           .write
		.ctrl_out_s1_readdata                                             (mm_interconnect_1_ctrl_out_s1_readdata),                                //                                                           .readdata
		.ctrl_out_s1_writedata                                            (mm_interconnect_1_ctrl_out_s1_writedata),                               //                                                           .writedata
		.ctrl_out_s1_chipselect                                           (mm_interconnect_1_ctrl_out_s1_chipselect),                              //                                                           .chipselect
		.dac_grad_spi_control_port_address                                (mm_interconnect_1_dac_grad_spi_control_port_address),                   //                                  dac_grad_spi_control_port.address
		.dac_grad_spi_control_port_write                                  (mm_interconnect_1_dac_grad_spi_control_port_write),                     //                                                           .write
		.dac_grad_spi_control_port_read                                   (mm_interconnect_1_dac_grad_spi_control_port_read),                      //                                                           .read
		.dac_grad_spi_control_port_readdata                               (mm_interconnect_1_dac_grad_spi_control_port_readdata),                  //                                                           .readdata
		.dac_grad_spi_control_port_writedata                              (mm_interconnect_1_dac_grad_spi_control_port_writedata),                 //                                                           .writedata
		.dac_grad_spi_control_port_chipselect                             (mm_interconnect_1_dac_grad_spi_control_port_chipselect),                //                                                           .chipselect
		.dconv_fifo_mem_in_csr_address                                    (mm_interconnect_1_dconv_fifo_mem_in_csr_address),                       //                                      dconv_fifo_mem_in_csr.address
		.dconv_fifo_mem_in_csr_write                                      (mm_interconnect_1_dconv_fifo_mem_in_csr_write),                         //                                                           .write
		.dconv_fifo_mem_in_csr_read                                       (mm_interconnect_1_dconv_fifo_mem_in_csr_read),                          //                                                           .read
		.dconv_fifo_mem_in_csr_readdata                                   (mm_interconnect_1_dconv_fifo_mem_in_csr_readdata),                      //                                                           .readdata
		.dconv_fifo_mem_in_csr_writedata                                  (mm_interconnect_1_dconv_fifo_mem_in_csr_writedata),                     //                                                           .writedata
		.dconv_fifo_mem_out_address                                       (mm_interconnect_1_dconv_fifo_mem_out_address),                          //                                         dconv_fifo_mem_out.address
		.dconv_fifo_mem_out_read                                          (mm_interconnect_1_dconv_fifo_mem_out_read),                             //                                                           .read
		.dconv_fifo_mem_out_readdata                                      (mm_interconnect_1_dconv_fifo_mem_out_readdata),                         //                                                           .readdata
		.dconv_fifo_mem_out_waitrequest                                   (mm_interconnect_1_dconv_fifo_mem_out_waitrequest),                      //                                                           .waitrequest
		.dconv_fifo_mem_q_in_csr_address                                  (mm_interconnect_1_dconv_fifo_mem_q_in_csr_address),                     //                                    dconv_fifo_mem_q_in_csr.address
		.dconv_fifo_mem_q_in_csr_write                                    (mm_interconnect_1_dconv_fifo_mem_q_in_csr_write),                       //                                                           .write
		.dconv_fifo_mem_q_in_csr_read                                     (mm_interconnect_1_dconv_fifo_mem_q_in_csr_read),                        //                                                           .read
		.dconv_fifo_mem_q_in_csr_readdata                                 (mm_interconnect_1_dconv_fifo_mem_q_in_csr_readdata),                    //                                                           .readdata
		.dconv_fifo_mem_q_in_csr_writedata                                (mm_interconnect_1_dconv_fifo_mem_q_in_csr_writedata),                   //                                                           .writedata
		.dconv_fifo_mem_q_out_address                                     (mm_interconnect_1_dconv_fifo_mem_q_out_address),                        //                                       dconv_fifo_mem_q_out.address
		.dconv_fifo_mem_q_out_read                                        (mm_interconnect_1_dconv_fifo_mem_q_out_read),                           //                                                           .read
		.dconv_fifo_mem_q_out_readdata                                    (mm_interconnect_1_dconv_fifo_mem_q_out_readdata),                       //                                                           .readdata
		.dconv_fifo_mem_q_out_waitrequest                                 (mm_interconnect_1_dconv_fifo_mem_q_out_waitrequest),                    //                                                           .waitrequest
		.dconv_fir_avalon_mm_slave_address                                (mm_interconnect_1_dconv_fir_avalon_mm_slave_address),                   //                                  dconv_fir_avalon_mm_slave.address
		.dconv_fir_avalon_mm_slave_write                                  (mm_interconnect_1_dconv_fir_avalon_mm_slave_write),                     //                                                           .write
		.dconv_fir_avalon_mm_slave_read                                   (mm_interconnect_1_dconv_fir_avalon_mm_slave_read),                      //                                                           .read
		.dconv_fir_avalon_mm_slave_readdata                               (mm_interconnect_1_dconv_fir_avalon_mm_slave_readdata),                  //                                                           .readdata
		.dconv_fir_avalon_mm_slave_writedata                              (mm_interconnect_1_dconv_fir_avalon_mm_slave_writedata),                 //                                                           .writedata
		.dconv_fir_avalon_mm_slave_readdatavalid                          (mm_interconnect_1_dconv_fir_avalon_mm_slave_readdatavalid),             //                                                           .readdatavalid
		.dconv_fir_q_avalon_mm_slave_address                              (mm_interconnect_1_dconv_fir_q_avalon_mm_slave_address),                 //                                dconv_fir_q_avalon_mm_slave.address
		.dconv_fir_q_avalon_mm_slave_write                                (mm_interconnect_1_dconv_fir_q_avalon_mm_slave_write),                   //                                                           .write
		.dconv_fir_q_avalon_mm_slave_read                                 (mm_interconnect_1_dconv_fir_q_avalon_mm_slave_read),                    //                                                           .read
		.dconv_fir_q_avalon_mm_slave_readdata                             (mm_interconnect_1_dconv_fir_q_avalon_mm_slave_readdata),                //                                                           .readdata
		.dconv_fir_q_avalon_mm_slave_writedata                            (mm_interconnect_1_dconv_fir_q_avalon_mm_slave_writedata),               //                                                           .writedata
		.dconv_fir_q_avalon_mm_slave_readdatavalid                        (mm_interconnect_1_dconv_fir_q_avalon_mm_slave_readdatavalid),           //                                                           .readdatavalid
		.dma_dconvi_control_port_slave_address                            (mm_interconnect_1_dma_dconvi_control_port_slave_address),               //                              dma_dconvi_control_port_slave.address
		.dma_dconvi_control_port_slave_write                              (mm_interconnect_1_dma_dconvi_control_port_slave_write),                 //                                                           .write
		.dma_dconvi_control_port_slave_readdata                           (mm_interconnect_1_dma_dconvi_control_port_slave_readdata),              //                                                           .readdata
		.dma_dconvi_control_port_slave_writedata                          (mm_interconnect_1_dma_dconvi_control_port_slave_writedata),             //                                                           .writedata
		.dma_dconvi_control_port_slave_chipselect                         (mm_interconnect_1_dma_dconvi_control_port_slave_chipselect),            //                                                           .chipselect
		.dma_dconvq_control_port_slave_address                            (mm_interconnect_1_dma_dconvq_control_port_slave_address),               //                              dma_dconvq_control_port_slave.address
		.dma_dconvq_control_port_slave_write                              (mm_interconnect_1_dma_dconvq_control_port_slave_write),                 //                                                           .write
		.dma_dconvq_control_port_slave_readdata                           (mm_interconnect_1_dma_dconvq_control_port_slave_readdata),              //                                                           .readdata
		.dma_dconvq_control_port_slave_writedata                          (mm_interconnect_1_dma_dconvq_control_port_slave_writedata),             //                                                           .writedata
		.dma_dconvq_control_port_slave_chipselect                         (mm_interconnect_1_dma_dconvq_control_port_slave_chipselect),            //                                                           .chipselect
		.dma_dummy_control_port_slave_address                             (mm_interconnect_1_dma_dummy_control_port_slave_address),                //                               dma_dummy_control_port_slave.address
		.dma_dummy_control_port_slave_write                               (mm_interconnect_1_dma_dummy_control_port_slave_write),                  //                                                           .write
		.dma_dummy_control_port_slave_readdata                            (mm_interconnect_1_dma_dummy_control_port_slave_readdata),               //                                                           .readdata
		.dma_dummy_control_port_slave_writedata                           (mm_interconnect_1_dma_dummy_control_port_slave_writedata),              //                                                           .writedata
		.dma_dummy_control_port_slave_chipselect                          (mm_interconnect_1_dma_dummy_control_port_slave_chipselect),             //                                                           .chipselect
		.dma_fifo_control_port_slave_address                              (mm_interconnect_1_dma_fifo_control_port_slave_address),                 //                                dma_fifo_control_port_slave.address
		.dma_fifo_control_port_slave_write                                (mm_interconnect_1_dma_fifo_control_port_slave_write),                   //                                                           .write
		.dma_fifo_control_port_slave_readdata                             (mm_interconnect_1_dma_fifo_control_port_slave_readdata),                //                                                           .readdata
		.dma_fifo_control_port_slave_writedata                            (mm_interconnect_1_dma_fifo_control_port_slave_writedata),               //                                                           .writedata
		.dma_fifo_control_port_slave_chipselect                           (mm_interconnect_1_dma_fifo_control_port_slave_chipselect),              //                                                           .chipselect
		.fifo_dummy_in_write                                              (mm_interconnect_1_fifo_dummy_in_write),                                 //                                              fifo_dummy_in.write
		.fifo_dummy_in_writedata                                          (mm_interconnect_1_fifo_dummy_in_writedata),                             //                                                           .writedata
		.fifo_dummy_in_waitrequest                                        (mm_interconnect_1_fifo_dummy_in_waitrequest),                           //                                                           .waitrequest
		.fifo_dummy_in_csr_address                                        (mm_interconnect_1_fifo_dummy_in_csr_address),                           //                                          fifo_dummy_in_csr.address
		.fifo_dummy_in_csr_write                                          (mm_interconnect_1_fifo_dummy_in_csr_write),                             //                                                           .write
		.fifo_dummy_in_csr_read                                           (mm_interconnect_1_fifo_dummy_in_csr_read),                              //                                                           .read
		.fifo_dummy_in_csr_readdata                                       (mm_interconnect_1_fifo_dummy_in_csr_readdata),                          //                                                           .readdata
		.fifo_dummy_in_csr_writedata                                      (mm_interconnect_1_fifo_dummy_in_csr_writedata),                         //                                                           .writedata
		.fifo_dummy_out_read                                              (mm_interconnect_1_fifo_dummy_out_read),                                 //                                             fifo_dummy_out.read
		.fifo_dummy_out_readdata                                          (mm_interconnect_1_fifo_dummy_out_readdata),                             //                                                           .readdata
		.fifo_dummy_out_waitrequest                                       (mm_interconnect_1_fifo_dummy_out_waitrequest),                          //                                                           .waitrequest
		.fifo_dummy64_in_in_address                                       (mm_interconnect_1_fifo_dummy64_in_in_address),                          //                                         fifo_dummy64_in_in.address
		.fifo_dummy64_in_in_write                                         (mm_interconnect_1_fifo_dummy64_in_in_write),                            //                                                           .write
		.fifo_dummy64_in_in_writedata                                     (mm_interconnect_1_fifo_dummy64_in_in_writedata),                        //                                                           .writedata
		.fifo_dummy64_in_in_waitrequest                                   (mm_interconnect_1_fifo_dummy64_in_in_waitrequest),                      //                                                           .waitrequest
		.fifo_dummy64_in_in_csr_address                                   (mm_interconnect_1_fifo_dummy64_in_in_csr_address),                      //                                     fifo_dummy64_in_in_csr.address
		.fifo_dummy64_in_in_csr_write                                     (mm_interconnect_1_fifo_dummy64_in_in_csr_write),                        //                                                           .write
		.fifo_dummy64_in_in_csr_read                                      (mm_interconnect_1_fifo_dummy64_in_in_csr_read),                         //                                                           .read
		.fifo_dummy64_in_in_csr_readdata                                  (mm_interconnect_1_fifo_dummy64_in_in_csr_readdata),                     //                                                           .readdata
		.fifo_dummy64_in_in_csr_writedata                                 (mm_interconnect_1_fifo_dummy64_in_in_csr_writedata),                    //                                                           .writedata
		.fifo_dummy64_out_in_csr_address                                  (mm_interconnect_1_fifo_dummy64_out_in_csr_address),                     //                                    fifo_dummy64_out_in_csr.address
		.fifo_dummy64_out_in_csr_write                                    (mm_interconnect_1_fifo_dummy64_out_in_csr_write),                       //                                                           .write
		.fifo_dummy64_out_in_csr_read                                     (mm_interconnect_1_fifo_dummy64_out_in_csr_read),                        //                                                           .read
		.fifo_dummy64_out_in_csr_readdata                                 (mm_interconnect_1_fifo_dummy64_out_in_csr_readdata),                    //                                                           .readdata
		.fifo_dummy64_out_in_csr_writedata                                (mm_interconnect_1_fifo_dummy64_out_in_csr_writedata),                   //                                                           .writedata
		.fifo_dummy64_out_out_address                                     (mm_interconnect_1_fifo_dummy64_out_out_address),                        //                                       fifo_dummy64_out_out.address
		.fifo_dummy64_out_out_read                                        (mm_interconnect_1_fifo_dummy64_out_out_read),                           //                                                           .read
		.fifo_dummy64_out_out_readdata                                    (mm_interconnect_1_fifo_dummy64_out_out_readdata),                       //                                                           .readdata
		.fifo_dummy64_out_out_waitrequest                                 (mm_interconnect_1_fifo_dummy64_out_out_waitrequest),                    //                                                           .waitrequest
		.i2c_ext_csr_address                                              (mm_interconnect_1_i2c_ext_csr_address),                                 //                                                i2c_ext_csr.address
		.i2c_ext_csr_write                                                (mm_interconnect_1_i2c_ext_csr_write),                                   //                                                           .write
		.i2c_ext_csr_read                                                 (mm_interconnect_1_i2c_ext_csr_read),                                    //                                                           .read
		.i2c_ext_csr_readdata                                             (mm_interconnect_1_i2c_ext_csr_readdata),                                //                                                           .readdata
		.i2c_ext_csr_writedata                                            (mm_interconnect_1_i2c_ext_csr_writedata),                               //                                                           .writedata
		.i2c_int_csr_address                                              (mm_interconnect_1_i2c_int_csr_address),                                 //                                                i2c_int_csr.address
		.i2c_int_csr_write                                                (mm_interconnect_1_i2c_int_csr_write),                                   //                                                           .write
		.i2c_int_csr_read                                                 (mm_interconnect_1_i2c_int_csr_read),                                    //                                                           .read
		.i2c_int_csr_readdata                                             (mm_interconnect_1_i2c_int_csr_readdata),                                //                                                           .readdata
		.i2c_int_csr_writedata                                            (mm_interconnect_1_i2c_int_csr_writedata),                               //                                                           .writedata
		.jtag_uart_avalon_jtag_slave_address                              (mm_interconnect_1_jtag_uart_avalon_jtag_slave_address),                 //                                jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                                (mm_interconnect_1_jtag_uart_avalon_jtag_slave_write),                   //                                                           .write
		.jtag_uart_avalon_jtag_slave_read                                 (mm_interconnect_1_jtag_uart_avalon_jtag_slave_read),                    //                                                           .read
		.jtag_uart_avalon_jtag_slave_readdata                             (mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata),                //                                                           .readdata
		.jtag_uart_avalon_jtag_slave_writedata                            (mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata),               //                                                           .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest                          (mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest),             //                                                           .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                           (mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect),              //                                                           .chipselect
		.nmr_parameters_adc_val_sub_s1_address                            (mm_interconnect_1_nmr_parameters_adc_val_sub_s1_address),               //                              nmr_parameters_adc_val_sub_s1.address
		.nmr_parameters_adc_val_sub_s1_write                              (mm_interconnect_1_nmr_parameters_adc_val_sub_s1_write),                 //                                                           .write
		.nmr_parameters_adc_val_sub_s1_readdata                           (mm_interconnect_1_nmr_parameters_adc_val_sub_s1_readdata),              //                                                           .readdata
		.nmr_parameters_adc_val_sub_s1_writedata                          (mm_interconnect_1_nmr_parameters_adc_val_sub_s1_writedata),             //                                                           .writedata
		.nmr_parameters_adc_val_sub_s1_chipselect                         (mm_interconnect_1_nmr_parameters_adc_val_sub_s1_chipselect),            //                                                           .chipselect
		.nmr_parameters_delay_nosig_s1_address                            (mm_interconnect_1_nmr_parameters_delay_nosig_s1_address),               //                              nmr_parameters_delay_nosig_s1.address
		.nmr_parameters_delay_nosig_s1_write                              (mm_interconnect_1_nmr_parameters_delay_nosig_s1_write),                 //                                                           .write
		.nmr_parameters_delay_nosig_s1_readdata                           (mm_interconnect_1_nmr_parameters_delay_nosig_s1_readdata),              //                                                           .readdata
		.nmr_parameters_delay_nosig_s1_writedata                          (mm_interconnect_1_nmr_parameters_delay_nosig_s1_writedata),             //                                                           .writedata
		.nmr_parameters_delay_nosig_s1_chipselect                         (mm_interconnect_1_nmr_parameters_delay_nosig_s1_chipselect),            //                                                           .chipselect
		.nmr_parameters_delay_sig_s1_address                              (mm_interconnect_1_nmr_parameters_delay_sig_s1_address),                 //                                nmr_parameters_delay_sig_s1.address
		.nmr_parameters_delay_sig_s1_write                                (mm_interconnect_1_nmr_parameters_delay_sig_s1_write),                   //                                                           .write
		.nmr_parameters_delay_sig_s1_readdata                             (mm_interconnect_1_nmr_parameters_delay_sig_s1_readdata),                //                                                           .readdata
		.nmr_parameters_delay_sig_s1_writedata                            (mm_interconnect_1_nmr_parameters_delay_sig_s1_writedata),               //                                                           .writedata
		.nmr_parameters_delay_sig_s1_chipselect                           (mm_interconnect_1_nmr_parameters_delay_sig_s1_chipselect),              //                                                           .chipselect
		.nmr_parameters_delay_t1_s1_address                               (mm_interconnect_1_nmr_parameters_delay_t1_s1_address),                  //                                 nmr_parameters_delay_t1_s1.address
		.nmr_parameters_delay_t1_s1_write                                 (mm_interconnect_1_nmr_parameters_delay_t1_s1_write),                    //                                                           .write
		.nmr_parameters_delay_t1_s1_readdata                              (mm_interconnect_1_nmr_parameters_delay_t1_s1_readdata),                 //                                                           .readdata
		.nmr_parameters_delay_t1_s1_writedata                             (mm_interconnect_1_nmr_parameters_delay_t1_s1_writedata),                //                                                           .writedata
		.nmr_parameters_delay_t1_s1_chipselect                            (mm_interconnect_1_nmr_parameters_delay_t1_s1_chipselect),               //                                                           .chipselect
		.nmr_parameters_echoes_per_scan_s1_address                        (mm_interconnect_1_nmr_parameters_echoes_per_scan_s1_address),           //                          nmr_parameters_echoes_per_scan_s1.address
		.nmr_parameters_echoes_per_scan_s1_write                          (mm_interconnect_1_nmr_parameters_echoes_per_scan_s1_write),             //                                                           .write
		.nmr_parameters_echoes_per_scan_s1_readdata                       (mm_interconnect_1_nmr_parameters_echoes_per_scan_s1_readdata),          //                                                           .readdata
		.nmr_parameters_echoes_per_scan_s1_writedata                      (mm_interconnect_1_nmr_parameters_echoes_per_scan_s1_writedata),         //                                                           .writedata
		.nmr_parameters_echoes_per_scan_s1_chipselect                     (mm_interconnect_1_nmr_parameters_echoes_per_scan_s1_chipselect),        //                                                           .chipselect
		.nmr_parameters_init_delay_s1_address                             (mm_interconnect_1_nmr_parameters_init_delay_s1_address),                //                               nmr_parameters_init_delay_s1.address
		.nmr_parameters_init_delay_s1_write                               (mm_interconnect_1_nmr_parameters_init_delay_s1_write),                  //                                                           .write
		.nmr_parameters_init_delay_s1_readdata                            (mm_interconnect_1_nmr_parameters_init_delay_s1_readdata),               //                                                           .readdata
		.nmr_parameters_init_delay_s1_writedata                           (mm_interconnect_1_nmr_parameters_init_delay_s1_writedata),              //                                                           .writedata
		.nmr_parameters_init_delay_s1_chipselect                          (mm_interconnect_1_nmr_parameters_init_delay_s1_chipselect),             //                                                           .chipselect
		.nmr_parameters_pulse_180deg_s1_address                           (mm_interconnect_1_nmr_parameters_pulse_180deg_s1_address),              //                             nmr_parameters_pulse_180deg_s1.address
		.nmr_parameters_pulse_180deg_s1_write                             (mm_interconnect_1_nmr_parameters_pulse_180deg_s1_write),                //                                                           .write
		.nmr_parameters_pulse_180deg_s1_readdata                          (mm_interconnect_1_nmr_parameters_pulse_180deg_s1_readdata),             //                                                           .readdata
		.nmr_parameters_pulse_180deg_s1_writedata                         (mm_interconnect_1_nmr_parameters_pulse_180deg_s1_writedata),            //                                                           .writedata
		.nmr_parameters_pulse_180deg_s1_chipselect                        (mm_interconnect_1_nmr_parameters_pulse_180deg_s1_chipselect),           //                                                           .chipselect
		.nmr_parameters_pulse_90deg_s1_address                            (mm_interconnect_1_nmr_parameters_pulse_90deg_s1_address),               //                              nmr_parameters_pulse_90deg_s1.address
		.nmr_parameters_pulse_90deg_s1_write                              (mm_interconnect_1_nmr_parameters_pulse_90deg_s1_write),                 //                                                           .write
		.nmr_parameters_pulse_90deg_s1_readdata                           (mm_interconnect_1_nmr_parameters_pulse_90deg_s1_readdata),              //                                                           .readdata
		.nmr_parameters_pulse_90deg_s1_writedata                          (mm_interconnect_1_nmr_parameters_pulse_90deg_s1_writedata),             //                                                           .writedata
		.nmr_parameters_pulse_90deg_s1_chipselect                         (mm_interconnect_1_nmr_parameters_pulse_90deg_s1_chipselect),            //                                                           .chipselect
		.nmr_parameters_pulse_t1_s1_address                               (mm_interconnect_1_nmr_parameters_pulse_t1_s1_address),                  //                                 nmr_parameters_pulse_t1_s1.address
		.nmr_parameters_pulse_t1_s1_write                                 (mm_interconnect_1_nmr_parameters_pulse_t1_s1_write),                    //                                                           .write
		.nmr_parameters_pulse_t1_s1_readdata                              (mm_interconnect_1_nmr_parameters_pulse_t1_s1_readdata),                 //                                                           .readdata
		.nmr_parameters_pulse_t1_s1_writedata                             (mm_interconnect_1_nmr_parameters_pulse_t1_s1_writedata),                //                                                           .writedata
		.nmr_parameters_pulse_t1_s1_chipselect                            (mm_interconnect_1_nmr_parameters_pulse_t1_s1_chipselect),               //                                                           .chipselect
		.nmr_parameters_rx_delay_s1_address                               (mm_interconnect_1_nmr_parameters_rx_delay_s1_address),                  //                                 nmr_parameters_rx_delay_s1.address
		.nmr_parameters_rx_delay_s1_write                                 (mm_interconnect_1_nmr_parameters_rx_delay_s1_write),                    //                                                           .write
		.nmr_parameters_rx_delay_s1_readdata                              (mm_interconnect_1_nmr_parameters_rx_delay_s1_readdata),                 //                                                           .readdata
		.nmr_parameters_rx_delay_s1_writedata                             (mm_interconnect_1_nmr_parameters_rx_delay_s1_writedata),                //                                                           .writedata
		.nmr_parameters_rx_delay_s1_chipselect                            (mm_interconnect_1_nmr_parameters_rx_delay_s1_chipselect),               //                                                           .chipselect
		.nmr_parameters_samples_per_echo_s1_address                       (mm_interconnect_1_nmr_parameters_samples_per_echo_s1_address),          //                         nmr_parameters_samples_per_echo_s1.address
		.nmr_parameters_samples_per_echo_s1_write                         (mm_interconnect_1_nmr_parameters_samples_per_echo_s1_write),            //                                                           .write
		.nmr_parameters_samples_per_echo_s1_readdata                      (mm_interconnect_1_nmr_parameters_samples_per_echo_s1_readdata),         //                                                           .readdata
		.nmr_parameters_samples_per_echo_s1_writedata                     (mm_interconnect_1_nmr_parameters_samples_per_echo_s1_writedata),        //                                                           .writedata
		.nmr_parameters_samples_per_echo_s1_chipselect                    (mm_interconnect_1_nmr_parameters_samples_per_echo_s1_chipselect),       //                                                           .chipselect
		.nmr_sys_pll_reconfig_mgmt_avalon_slave_address                   (mm_interconnect_1_nmr_sys_pll_reconfig_mgmt_avalon_slave_address),      //                     nmr_sys_pll_reconfig_mgmt_avalon_slave.address
		.nmr_sys_pll_reconfig_mgmt_avalon_slave_write                     (mm_interconnect_1_nmr_sys_pll_reconfig_mgmt_avalon_slave_write),        //                                                           .write
		.nmr_sys_pll_reconfig_mgmt_avalon_slave_read                      (mm_interconnect_1_nmr_sys_pll_reconfig_mgmt_avalon_slave_read),         //                                                           .read
		.nmr_sys_pll_reconfig_mgmt_avalon_slave_readdata                  (mm_interconnect_1_nmr_sys_pll_reconfig_mgmt_avalon_slave_readdata),     //                                                           .readdata
		.nmr_sys_pll_reconfig_mgmt_avalon_slave_writedata                 (mm_interconnect_1_nmr_sys_pll_reconfig_mgmt_avalon_slave_writedata),    //                                                           .writedata
		.nmr_sys_pll_reconfig_mgmt_avalon_slave_waitrequest               (mm_interconnect_1_nmr_sys_pll_reconfig_mgmt_avalon_slave_waitrequest),  //                                                           .waitrequest
		.sdram_s1_address                                                 (mm_interconnect_1_sdram_s1_address),                                    //                                                   sdram_s1.address
		.sdram_s1_write                                                   (mm_interconnect_1_sdram_s1_write),                                      //                                                           .write
		.sdram_s1_read                                                    (mm_interconnect_1_sdram_s1_read),                                       //                                                           .read
		.sdram_s1_readdata                                                (mm_interconnect_1_sdram_s1_readdata),                                   //                                                           .readdata
		.sdram_s1_writedata                                               (mm_interconnect_1_sdram_s1_writedata),                                  //                                                           .writedata
		.sdram_s1_byteenable                                              (mm_interconnect_1_sdram_s1_byteenable),                                 //                                                           .byteenable
		.sdram_s1_readdatavalid                                           (mm_interconnect_1_sdram_s1_readdatavalid),                              //                                                           .readdatavalid
		.sdram_s1_waitrequest                                             (mm_interconnect_1_sdram_s1_waitrequest),                                //                                                           .waitrequest
		.sdram_s1_chipselect                                              (mm_interconnect_1_sdram_s1_chipselect),                                 //                                                           .chipselect
		.spi_afe_relays_spi_control_port_address                          (mm_interconnect_1_spi_afe_relays_spi_control_port_address),             //                            spi_afe_relays_spi_control_port.address
		.spi_afe_relays_spi_control_port_write                            (mm_interconnect_1_spi_afe_relays_spi_control_port_write),               //                                                           .write
		.spi_afe_relays_spi_control_port_read                             (mm_interconnect_1_spi_afe_relays_spi_control_port_read),                //                                                           .read
		.spi_afe_relays_spi_control_port_readdata                         (mm_interconnect_1_spi_afe_relays_spi_control_port_readdata),            //                                                           .readdata
		.spi_afe_relays_spi_control_port_writedata                        (mm_interconnect_1_spi_afe_relays_spi_control_port_writedata),           //                                                           .writedata
		.spi_afe_relays_spi_control_port_chipselect                       (mm_interconnect_1_spi_afe_relays_spi_control_port_chipselect),          //                                                           .chipselect
		.spi_mtch_ntwrk_spi_control_port_address                          (mm_interconnect_1_spi_mtch_ntwrk_spi_control_port_address),             //                            spi_mtch_ntwrk_spi_control_port.address
		.spi_mtch_ntwrk_spi_control_port_write                            (mm_interconnect_1_spi_mtch_ntwrk_spi_control_port_write),               //                                                           .write
		.spi_mtch_ntwrk_spi_control_port_read                             (mm_interconnect_1_spi_mtch_ntwrk_spi_control_port_read),                //                                                           .read
		.spi_mtch_ntwrk_spi_control_port_readdata                         (mm_interconnect_1_spi_mtch_ntwrk_spi_control_port_readdata),            //                                                           .readdata
		.spi_mtch_ntwrk_spi_control_port_writedata                        (mm_interconnect_1_spi_mtch_ntwrk_spi_control_port_writedata),           //                                                           .writedata
		.spi_mtch_ntwrk_spi_control_port_chipselect                       (mm_interconnect_1_spi_mtch_ntwrk_spi_control_port_chipselect),          //                                                           .chipselect
		.switches_s1_address                                              (mm_interconnect_1_switches_s1_address),                                 //                                                switches_s1.address
		.switches_s1_readdata                                             (mm_interconnect_1_switches_s1_readdata),                                //                                                           .readdata
		.sysid_qsys_control_slave_address                                 (mm_interconnect_1_sysid_qsys_control_slave_address),                    //                                   sysid_qsys_control_slave.address
		.sysid_qsys_control_slave_readdata                                (mm_interconnect_1_sysid_qsys_control_slave_readdata)                    //                                                           .readdata
	);

	soc_system_v5_irq_mapper irq_mapper (
		.clk           (),                         //       clk.clk
		.reset         (),                         // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq), // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq), // receiver1.irq
		.sender_irq    (hps_0_f2h_irq0_irq)        //    sender.irq
	);

	soc_system_v5_irq_mapper_001 irq_mapper_001 (
		.clk           (),                             //       clk.clk
		.reset         (),                             // clk_reset.reset
		.receiver0_irq (irq_mapper_001_receiver0_irq), // receiver0.irq
		.receiver1_irq (irq_mapper_001_receiver1_irq), // receiver1.irq
		.receiver2_irq (irq_mapper_001_receiver2_irq), // receiver2.irq
		.receiver3_irq (irq_mapper_001_receiver3_irq), // receiver3.irq
		.receiver4_irq (irq_mapper_001_receiver4_irq), // receiver4.irq
		.receiver5_irq (irq_mapper_001_receiver5_irq), // receiver5.irq
		.receiver6_irq (irq_mapper_001_receiver6_irq), // receiver6.irq
		.receiver7_irq (irq_mapper_001_receiver7_irq), // receiver7.irq
		.sender_irq    (hps_0_f2h_irq1_irq)            //    sender.irq
	);

	soc_system_v5_avalon_st_adapter #(
		.inBitsPerSymbol (16),
		.inUsePackets    (0),
		.inDataWidth     (16),
		.inChannelWidth  (0),
		.inErrorWidth    (0),
		.inUseEmptyPort  (0),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (32),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (0),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (1)
	) avalon_st_adapter (
		.in_clk_0_clk   (clk_clk),                            // in_clk_0.clk
		.in_rst_0_reset (rst_controller_001_reset_out_reset), // in_rst_0.reset
		.in_0_data      (adc_fifo_dc_out_data),               //     in_0.data
		.in_0_valid     (adc_fifo_dc_out_valid),              //         .valid
		.in_0_ready     (adc_fifo_dc_out_ready),              //         .ready
		.out_0_data     (avalon_st_adapter_out_0_data),       //    out_0.data
		.out_0_valid    (avalon_st_adapter_out_0_valid),      //         .valid
		.out_0_ready    (avalon_st_adapter_out_0_ready)       //         .ready
	);

	soc_system_v5_avalon_st_adapter_001 #(
		.inBitsPerSymbol (32),
		.inUsePackets    (0),
		.inDataWidth     (32),
		.inChannelWidth  (0),
		.inErrorWidth    (0),
		.inUseEmptyPort  (0),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (32),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (0),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (1)
	) avalon_st_adapter_001 (
		.in_clk_0_clk   (clk_clk),                            // in_clk_0.clk
		.in_rst_0_reset (rst_controller_001_reset_out_reset), // in_rst_0.reset
		.in_0_data      (dconv_fifo_dc_out_data),             //     in_0.data
		.in_0_valid     (dconv_fifo_dc_out_valid),            //         .valid
		.in_0_ready     (dconv_fifo_dc_out_ready),            //         .ready
		.out_0_data     (avalon_st_adapter_001_out_0_data),   //    out_0.data
		.out_0_valid    (avalon_st_adapter_001_out_0_valid),  //         .valid
		.out_0_ready    (avalon_st_adapter_001_out_0_ready)   //         .ready
	);

	soc_system_v5_avalon_st_adapter_001 #(
		.inBitsPerSymbol (32),
		.inUsePackets    (0),
		.inDataWidth     (32),
		.inChannelWidth  (0),
		.inErrorWidth    (0),
		.inUseEmptyPort  (0),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (32),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (0),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (1)
	) avalon_st_adapter_002 (
		.in_clk_0_clk   (clk_clk),                            // in_clk_0.clk
		.in_rst_0_reset (rst_controller_001_reset_out_reset), // in_rst_0.reset
		.in_0_data      (dconv_fifo_dc_q_out_data),           //     in_0.data
		.in_0_valid     (dconv_fifo_dc_q_out_valid),          //         .valid
		.in_0_ready     (dconv_fifo_dc_q_out_ready),          //         .ready
		.out_0_data     (avalon_st_adapter_002_out_0_data),   //    out_0.data
		.out_0_valid    (avalon_st_adapter_002_out_0_valid),  //         .valid
		.out_0_ready    (avalon_st_adapter_002_out_0_ready)   //         .ready
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.reset_in1      (fifo_rst_reset),                 // reset_in1.reset
		.clk            (fifo_clk_bridge_in_clk),         //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (fifo_rst_reset),                     // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (gp_pll_outclk0_clk),                 //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_004 (
		.reset_in0      (~hps_0_h2f_reset_reset_n),           // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_004_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
