-- soc_system_v5_dconv_fifo_dc.vhd

-- Generated using ACDS version 17.1 590

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity soc_system_v5_dconv_fifo_dc is
	generic (
		SYMBOLS_PER_BEAT   : integer := 1;
		BITS_PER_SYMBOL    : integer := 32;
		FIFO_DEPTH         : integer := 32768;
		CHANNEL_WIDTH      : integer := 0;
		ERROR_WIDTH        : integer := 0;
		USE_PACKETS        : integer := 0;
		USE_IN_FILL_LEVEL  : integer := 0;
		USE_OUT_FILL_LEVEL : integer := 0;
		WR_SYNC_DEPTH      : integer := 3;
		RD_SYNC_DEPTH      : integer := 3
	);
	port (
		in_clk            : in  std_logic                     := '0';             --        in_clk.clk
		in_reset_n        : in  std_logic                     := '0';             --  in_clk_reset.reset_n
		out_clk           : in  std_logic                     := '0';             --       out_clk.clk
		out_reset_n       : in  std_logic                     := '0';             -- out_clk_reset.reset_n
		in_data           : in  std_logic_vector(31 downto 0) := (others => '0'); --            in.data
		in_valid          : in  std_logic                     := '0';             --              .valid
		in_ready          : out std_logic;                                        --              .ready
		out_data          : out std_logic_vector(31 downto 0);                    --           out.data
		out_valid         : out std_logic;                                        --              .valid
		out_ready         : in  std_logic                     := '0';             --              .ready
		in_channel        : in  std_logic_vector(0 downto 0)  := (others => '0');
		in_csr_address    : in  std_logic                     := '0';
		in_csr_read       : in  std_logic                     := '0';
		in_csr_readdata   : out std_logic_vector(31 downto 0);
		in_csr_write      : in  std_logic                     := '0';
		in_csr_writedata  : in  std_logic_vector(31 downto 0) := (others => '0');
		in_empty          : in  std_logic_vector(0 downto 0)  := (others => '0');
		in_endofpacket    : in  std_logic                     := '0';
		in_error          : in  std_logic_vector(0 downto 0)  := (others => '0');
		in_startofpacket  : in  std_logic                     := '0';
		out_channel       : out std_logic_vector(0 downto 0);
		out_csr_address   : in  std_logic                     := '0';
		out_csr_read      : in  std_logic                     := '0';
		out_csr_readdata  : out std_logic_vector(31 downto 0);
		out_csr_write     : in  std_logic                     := '0';
		out_csr_writedata : in  std_logic_vector(31 downto 0) := (others => '0');
		out_empty         : out std_logic_vector(0 downto 0);
		out_endofpacket   : out std_logic;
		out_error         : out std_logic_vector(0 downto 0);
		out_startofpacket : out std_logic;
		space_avail_data  : out std_logic_vector(15 downto 0)
	);
end entity soc_system_v5_dconv_fifo_dc;

architecture rtl of soc_system_v5_dconv_fifo_dc is
	component altera_avalon_dc_fifo is
		generic (
			SYMBOLS_PER_BEAT   : integer := 1;
			BITS_PER_SYMBOL    : integer := 8;
			FIFO_DEPTH         : integer := 16;
			CHANNEL_WIDTH      : integer := 0;
			ERROR_WIDTH        : integer := 0;
			USE_PACKETS        : integer := 0;
			USE_IN_FILL_LEVEL  : integer := 0;
			USE_OUT_FILL_LEVEL : integer := 0;
			WR_SYNC_DEPTH      : integer := 3;
			RD_SYNC_DEPTH      : integer := 3
		);
		port (
			in_clk            : in  std_logic                     := 'X';             -- clk
			in_reset_n        : in  std_logic                     := 'X';             -- reset_n
			out_clk           : in  std_logic                     := 'X';             -- clk
			out_reset_n       : in  std_logic                     := 'X';             -- reset_n
			in_data           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			in_valid          : in  std_logic                     := 'X';             -- valid
			in_ready          : out std_logic;                                        -- ready
			out_data          : out std_logic_vector(31 downto 0);                    -- data
			out_valid         : out std_logic;                                        -- valid
			out_ready         : in  std_logic                     := 'X';             -- ready
			in_csr_address    : in  std_logic                     := 'X';             -- address
			in_csr_read       : in  std_logic                     := 'X';             -- read
			in_csr_write      : in  std_logic                     := 'X';             -- write
			in_csr_readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_csr_writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			out_csr_address   : in  std_logic                     := 'X';             -- address
			out_csr_read      : in  std_logic                     := 'X';             -- read
			out_csr_write     : in  std_logic                     := 'X';             -- write
			out_csr_readdata  : out std_logic_vector(31 downto 0);                    -- readdata
			out_csr_writedata : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			out_startofpacket : out std_logic;                                        -- startofpacket
			out_endofpacket   : out std_logic;                                        -- endofpacket
			in_empty          : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- empty
			out_empty         : out std_logic_vector(0 downto 0);                     -- empty
			in_error          : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- error
			out_error         : out std_logic_vector(0 downto 0);                     -- error
			in_channel        : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- channel
			out_channel       : out std_logic_vector(0 downto 0);                     -- channel
			space_avail_data  : out std_logic_vector(15 downto 0)                     -- data
		);
	end component altera_avalon_dc_fifo;

begin

	dconv_fifo_dc : component altera_avalon_dc_fifo
		generic map (
			SYMBOLS_PER_BEAT   => SYMBOLS_PER_BEAT,
			BITS_PER_SYMBOL    => BITS_PER_SYMBOL,
			FIFO_DEPTH         => FIFO_DEPTH,
			CHANNEL_WIDTH      => CHANNEL_WIDTH,
			ERROR_WIDTH        => ERROR_WIDTH,
			USE_PACKETS        => USE_PACKETS,
			USE_IN_FILL_LEVEL  => USE_IN_FILL_LEVEL,
			USE_OUT_FILL_LEVEL => USE_OUT_FILL_LEVEL,
			WR_SYNC_DEPTH      => WR_SYNC_DEPTH,
			RD_SYNC_DEPTH      => RD_SYNC_DEPTH
		)
		port map (
			in_clk            => in_clk,                             --        in_clk.clk
			in_reset_n        => in_reset_n,                         --  in_clk_reset.reset_n
			out_clk           => out_clk,                            --       out_clk.clk
			out_reset_n       => out_reset_n,                        -- out_clk_reset.reset_n
			in_data           => in_data,                            --            in.data
			in_valid          => in_valid,                           --              .valid
			in_ready          => in_ready,                           --              .ready
			out_data          => out_data,                           --           out.data
			out_valid         => out_valid,                          --              .valid
			out_ready         => out_ready,                          --              .ready
			in_csr_address    => '0',                                --   (terminated)
			in_csr_read       => '0',                                --   (terminated)
			in_csr_write      => '0',                                --   (terminated)
			in_csr_readdata   => open,                               --   (terminated)
			in_csr_writedata  => "00000000000000000000000000000000", --   (terminated)
			out_csr_address   => '0',                                --   (terminated)
			out_csr_read      => '0',                                --   (terminated)
			out_csr_write     => '0',                                --   (terminated)
			out_csr_readdata  => open,                               --   (terminated)
			out_csr_writedata => "00000000000000000000000000000000", --   (terminated)
			in_startofpacket  => '0',                                --   (terminated)
			in_endofpacket    => '0',                                --   (terminated)
			out_startofpacket => open,                               --   (terminated)
			out_endofpacket   => open,                               --   (terminated)
			in_empty          => "0",                                --   (terminated)
			out_empty         => open,                               --   (terminated)
			in_error          => "0",                                --   (terminated)
			out_error         => open,                               --   (terminated)
			in_channel        => "0",                                --   (terminated)
			out_channel       => open,                               --   (terminated)
			space_avail_data  => open                                --   (terminated)
		);

end architecture rtl; -- of soc_system_v5_dconv_fifo_dc
