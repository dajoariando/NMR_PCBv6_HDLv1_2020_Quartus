-- soc_system_v5_nmr_parameters.vhd

-- Generated using ACDS version 17.1 590

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity soc_system_v5_nmr_parameters is
	port (
		adc_val_sub_clk_clk                         : in  std_logic                     := '0';             --                      adc_val_sub_clk.clk
		adc_val_sub_external_connection_export      : out std_logic_vector(31 downto 0);                    --      adc_val_sub_external_connection.export
		adc_val_sub_reset_reset_n                   : in  std_logic                     := '0';             --                    adc_val_sub_reset.reset_n
		adc_val_sub_s1_address                      : in  std_logic_vector(1 downto 0)  := (others => '0'); --                       adc_val_sub_s1.address
		adc_val_sub_s1_write_n                      : in  std_logic                     := '0';             --                                     .write_n
		adc_val_sub_s1_writedata                    : in  std_logic_vector(31 downto 0) := (others => '0'); --                                     .writedata
		adc_val_sub_s1_chipselect                   : in  std_logic                     := '0';             --                                     .chipselect
		adc_val_sub_s1_readdata                     : out std_logic_vector(31 downto 0);                    --                                     .readdata
		delay_nosig_clk_clk                         : in  std_logic                     := '0';             --                      delay_nosig_clk.clk
		delay_nosig_external_connection_export      : out std_logic_vector(31 downto 0);                    --      delay_nosig_external_connection.export
		delay_nosig_reset_reset_n                   : in  std_logic                     := '0';             --                    delay_nosig_reset.reset_n
		delay_nosig_s1_address                      : in  std_logic_vector(1 downto 0)  := (others => '0'); --                       delay_nosig_s1.address
		delay_nosig_s1_write_n                      : in  std_logic                     := '0';             --                                     .write_n
		delay_nosig_s1_writedata                    : in  std_logic_vector(31 downto 0) := (others => '0'); --                                     .writedata
		delay_nosig_s1_chipselect                   : in  std_logic                     := '0';             --                                     .chipselect
		delay_nosig_s1_readdata                     : out std_logic_vector(31 downto 0);                    --                                     .readdata
		delay_sig_clk_clk                           : in  std_logic                     := '0';             --                        delay_sig_clk.clk
		delay_sig_external_connection_export        : out std_logic_vector(31 downto 0);                    --        delay_sig_external_connection.export
		delay_sig_reset_reset_n                     : in  std_logic                     := '0';             --                      delay_sig_reset.reset_n
		delay_sig_s1_address                        : in  std_logic_vector(1 downto 0)  := (others => '0'); --                         delay_sig_s1.address
		delay_sig_s1_write_n                        : in  std_logic                     := '0';             --                                     .write_n
		delay_sig_s1_writedata                      : in  std_logic_vector(31 downto 0) := (others => '0'); --                                     .writedata
		delay_sig_s1_chipselect                     : in  std_logic                     := '0';             --                                     .chipselect
		delay_sig_s1_readdata                       : out std_logic_vector(31 downto 0);                    --                                     .readdata
		delay_t1_clk_clk                            : in  std_logic                     := '0';             --                         delay_t1_clk.clk
		delay_t1_external_connection_export         : out std_logic_vector(31 downto 0);                    --         delay_t1_external_connection.export
		delay_t1_reset_reset_n                      : in  std_logic                     := '0';             --                       delay_t1_reset.reset_n
		delay_t1_s1_address                         : in  std_logic_vector(1 downto 0)  := (others => '0'); --                          delay_t1_s1.address
		delay_t1_s1_write_n                         : in  std_logic                     := '0';             --                                     .write_n
		delay_t1_s1_writedata                       : in  std_logic_vector(31 downto 0) := (others => '0'); --                                     .writedata
		delay_t1_s1_chipselect                      : in  std_logic                     := '0';             --                                     .chipselect
		delay_t1_s1_readdata                        : out std_logic_vector(31 downto 0);                    --                                     .readdata
		echoes_per_scan_clk_clk                     : in  std_logic                     := '0';             --                  echoes_per_scan_clk.clk
		echoes_per_scan_external_connection_export  : out std_logic_vector(31 downto 0);                    --  echoes_per_scan_external_connection.export
		echoes_per_scan_reset_reset_n               : in  std_logic                     := '0';             --                echoes_per_scan_reset.reset_n
		echoes_per_scan_s1_address                  : in  std_logic_vector(1 downto 0)  := (others => '0'); --                   echoes_per_scan_s1.address
		echoes_per_scan_s1_write_n                  : in  std_logic                     := '0';             --                                     .write_n
		echoes_per_scan_s1_writedata                : in  std_logic_vector(31 downto 0) := (others => '0'); --                                     .writedata
		echoes_per_scan_s1_chipselect               : in  std_logic                     := '0';             --                                     .chipselect
		echoes_per_scan_s1_readdata                 : out std_logic_vector(31 downto 0);                    --                                     .readdata
		init_delay_clk_clk                          : in  std_logic                     := '0';             --                       init_delay_clk.clk
		init_delay_external_connection_export       : out std_logic_vector(31 downto 0);                    --       init_delay_external_connection.export
		init_delay_reset_reset_n                    : in  std_logic                     := '0';             --                     init_delay_reset.reset_n
		init_delay_s1_address                       : in  std_logic_vector(1 downto 0)  := (others => '0'); --                        init_delay_s1.address
		init_delay_s1_write_n                       : in  std_logic                     := '0';             --                                     .write_n
		init_delay_s1_writedata                     : in  std_logic_vector(31 downto 0) := (others => '0'); --                                     .writedata
		init_delay_s1_chipselect                    : in  std_logic                     := '0';             --                                     .chipselect
		init_delay_s1_readdata                      : out std_logic_vector(31 downto 0);                    --                                     .readdata
		pulse_180deg_clk_clk                        : in  std_logic                     := '0';             --                     pulse_180deg_clk.clk
		pulse_180deg_external_connection_export     : out std_logic_vector(31 downto 0);                    --     pulse_180deg_external_connection.export
		pulse_180deg_reset_reset_n                  : in  std_logic                     := '0';             --                   pulse_180deg_reset.reset_n
		pulse_180deg_s1_address                     : in  std_logic_vector(1 downto 0)  := (others => '0'); --                      pulse_180deg_s1.address
		pulse_180deg_s1_write_n                     : in  std_logic                     := '0';             --                                     .write_n
		pulse_180deg_s1_writedata                   : in  std_logic_vector(31 downto 0) := (others => '0'); --                                     .writedata
		pulse_180deg_s1_chipselect                  : in  std_logic                     := '0';             --                                     .chipselect
		pulse_180deg_s1_readdata                    : out std_logic_vector(31 downto 0);                    --                                     .readdata
		pulse_90deg_clk_clk                         : in  std_logic                     := '0';             --                      pulse_90deg_clk.clk
		pulse_90deg_external_connection_export      : out std_logic_vector(31 downto 0);                    --      pulse_90deg_external_connection.export
		pulse_90deg_reset_reset_n                   : in  std_logic                     := '0';             --                    pulse_90deg_reset.reset_n
		pulse_90deg_s1_address                      : in  std_logic_vector(1 downto 0)  := (others => '0'); --                       pulse_90deg_s1.address
		pulse_90deg_s1_write_n                      : in  std_logic                     := '0';             --                                     .write_n
		pulse_90deg_s1_writedata                    : in  std_logic_vector(31 downto 0) := (others => '0'); --                                     .writedata
		pulse_90deg_s1_chipselect                   : in  std_logic                     := '0';             --                                     .chipselect
		pulse_90deg_s1_readdata                     : out std_logic_vector(31 downto 0);                    --                                     .readdata
		pulse_t1_clk_clk                            : in  std_logic                     := '0';             --                         pulse_t1_clk.clk
		pulse_t1_external_connection_export         : out std_logic_vector(31 downto 0);                    --         pulse_t1_external_connection.export
		pulse_t1_reset_reset_n                      : in  std_logic                     := '0';             --                       pulse_t1_reset.reset_n
		pulse_t1_s1_address                         : in  std_logic_vector(1 downto 0)  := (others => '0'); --                          pulse_t1_s1.address
		pulse_t1_s1_write_n                         : in  std_logic                     := '0';             --                                     .write_n
		pulse_t1_s1_writedata                       : in  std_logic_vector(31 downto 0) := (others => '0'); --                                     .writedata
		pulse_t1_s1_chipselect                      : in  std_logic                     := '0';             --                                     .chipselect
		pulse_t1_s1_readdata                        : out std_logic_vector(31 downto 0);                    --                                     .readdata
		rx_delay_clk_clk                            : in  std_logic                     := '0';             --                         rx_delay_clk.clk
		rx_delay_external_connection_export         : out std_logic_vector(31 downto 0);                    --         rx_delay_external_connection.export
		rx_delay_reset_reset_n                      : in  std_logic                     := '0';             --                       rx_delay_reset.reset_n
		rx_delay_s1_address                         : in  std_logic_vector(1 downto 0)  := (others => '0'); --                          rx_delay_s1.address
		rx_delay_s1_write_n                         : in  std_logic                     := '0';             --                                     .write_n
		rx_delay_s1_writedata                       : in  std_logic_vector(31 downto 0) := (others => '0'); --                                     .writedata
		rx_delay_s1_chipselect                      : in  std_logic                     := '0';             --                                     .chipselect
		rx_delay_s1_readdata                        : out std_logic_vector(31 downto 0);                    --                                     .readdata
		samples_per_echo_clk_clk                    : in  std_logic                     := '0';             --                 samples_per_echo_clk.clk
		samples_per_echo_external_connection_export : out std_logic_vector(31 downto 0);                    -- samples_per_echo_external_connection.export
		samples_per_echo_reset_reset_n              : in  std_logic                     := '0';             --               samples_per_echo_reset.reset_n
		samples_per_echo_s1_address                 : in  std_logic_vector(1 downto 0)  := (others => '0'); --                  samples_per_echo_s1.address
		samples_per_echo_s1_write_n                 : in  std_logic                     := '0';             --                                     .write_n
		samples_per_echo_s1_writedata               : in  std_logic_vector(31 downto 0) := (others => '0'); --                                     .writedata
		samples_per_echo_s1_chipselect              : in  std_logic                     := '0';             --                                     .chipselect
		samples_per_echo_s1_readdata                : out std_logic_vector(31 downto 0)                     --                                     .readdata
	);
end entity soc_system_v5_nmr_parameters;

architecture rtl of soc_system_v5_nmr_parameters is
	component soc_system_v5_nmr_parameters_adc_val_sub is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(31 downto 0)                     -- export
		);
	end component soc_system_v5_nmr_parameters_adc_val_sub;

	component soc_system_v5_nmr_parameters_delay_nosig is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(31 downto 0)                     -- export
		);
	end component soc_system_v5_nmr_parameters_delay_nosig;

	component soc_system_v5_nmr_parameters_delay_t1 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(31 downto 0)                     -- export
		);
	end component soc_system_v5_nmr_parameters_delay_t1;

	component soc_system_v5_nmr_parameters_samples_per_echo is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(31 downto 0)                     -- export
		);
	end component soc_system_v5_nmr_parameters_samples_per_echo;

begin

	adc_val_sub : component soc_system_v5_nmr_parameters_adc_val_sub
		port map (
			clk        => adc_val_sub_clk_clk,                    --                 clk.clk
			reset_n    => adc_val_sub_reset_reset_n,              --               reset.reset_n
			address    => adc_val_sub_s1_address,                 --                  s1.address
			write_n    => adc_val_sub_s1_write_n,                 --                    .write_n
			writedata  => adc_val_sub_s1_writedata,               --                    .writedata
			chipselect => adc_val_sub_s1_chipselect,              --                    .chipselect
			readdata   => adc_val_sub_s1_readdata,                --                    .readdata
			out_port   => adc_val_sub_external_connection_export  -- external_connection.export
		);

	delay_nosig : component soc_system_v5_nmr_parameters_delay_nosig
		port map (
			clk        => delay_nosig_clk_clk,                    --                 clk.clk
			reset_n    => delay_nosig_reset_reset_n,              --               reset.reset_n
			address    => delay_nosig_s1_address,                 --                  s1.address
			write_n    => delay_nosig_s1_write_n,                 --                    .write_n
			writedata  => delay_nosig_s1_writedata,               --                    .writedata
			chipselect => delay_nosig_s1_chipselect,              --                    .chipselect
			readdata   => delay_nosig_s1_readdata,                --                    .readdata
			out_port   => delay_nosig_external_connection_export  -- external_connection.export
		);

	delay_sig : component soc_system_v5_nmr_parameters_delay_nosig
		port map (
			clk        => delay_sig_clk_clk,                    --                 clk.clk
			reset_n    => delay_sig_reset_reset_n,              --               reset.reset_n
			address    => delay_sig_s1_address,                 --                  s1.address
			write_n    => delay_sig_s1_write_n,                 --                    .write_n
			writedata  => delay_sig_s1_writedata,               --                    .writedata
			chipselect => delay_sig_s1_chipselect,              --                    .chipselect
			readdata   => delay_sig_s1_readdata,                --                    .readdata
			out_port   => delay_sig_external_connection_export  -- external_connection.export
		);

	delay_t1 : component soc_system_v5_nmr_parameters_delay_t1
		port map (
			clk        => delay_t1_clk_clk,                    --                 clk.clk
			reset_n    => delay_t1_reset_reset_n,              --               reset.reset_n
			address    => delay_t1_s1_address,                 --                  s1.address
			write_n    => delay_t1_s1_write_n,                 --                    .write_n
			writedata  => delay_t1_s1_writedata,               --                    .writedata
			chipselect => delay_t1_s1_chipselect,              --                    .chipselect
			readdata   => delay_t1_s1_readdata,                --                    .readdata
			out_port   => delay_t1_external_connection_export  -- external_connection.export
		);

	echoes_per_scan : component soc_system_v5_nmr_parameters_delay_t1
		port map (
			clk        => echoes_per_scan_clk_clk,                    --                 clk.clk
			reset_n    => echoes_per_scan_reset_reset_n,              --               reset.reset_n
			address    => echoes_per_scan_s1_address,                 --                  s1.address
			write_n    => echoes_per_scan_s1_write_n,                 --                    .write_n
			writedata  => echoes_per_scan_s1_writedata,               --                    .writedata
			chipselect => echoes_per_scan_s1_chipselect,              --                    .chipselect
			readdata   => echoes_per_scan_s1_readdata,                --                    .readdata
			out_port   => echoes_per_scan_external_connection_export  -- external_connection.export
		);

	init_delay : component soc_system_v5_nmr_parameters_delay_t1
		port map (
			clk        => init_delay_clk_clk,                    --                 clk.clk
			reset_n    => init_delay_reset_reset_n,              --               reset.reset_n
			address    => init_delay_s1_address,                 --                  s1.address
			write_n    => init_delay_s1_write_n,                 --                    .write_n
			writedata  => init_delay_s1_writedata,               --                    .writedata
			chipselect => init_delay_s1_chipselect,              --                    .chipselect
			readdata   => init_delay_s1_readdata,                --                    .readdata
			out_port   => init_delay_external_connection_export  -- external_connection.export
		);

	pulse_180deg : component soc_system_v5_nmr_parameters_delay_nosig
		port map (
			clk        => pulse_180deg_clk_clk,                    --                 clk.clk
			reset_n    => pulse_180deg_reset_reset_n,              --               reset.reset_n
			address    => pulse_180deg_s1_address,                 --                  s1.address
			write_n    => pulse_180deg_s1_write_n,                 --                    .write_n
			writedata  => pulse_180deg_s1_writedata,               --                    .writedata
			chipselect => pulse_180deg_s1_chipselect,              --                    .chipselect
			readdata   => pulse_180deg_s1_readdata,                --                    .readdata
			out_port   => pulse_180deg_external_connection_export  -- external_connection.export
		);

	pulse_90deg : component soc_system_v5_nmr_parameters_delay_nosig
		port map (
			clk        => pulse_90deg_clk_clk,                    --                 clk.clk
			reset_n    => pulse_90deg_reset_reset_n,              --               reset.reset_n
			address    => pulse_90deg_s1_address,                 --                  s1.address
			write_n    => pulse_90deg_s1_write_n,                 --                    .write_n
			writedata  => pulse_90deg_s1_writedata,               --                    .writedata
			chipselect => pulse_90deg_s1_chipselect,              --                    .chipselect
			readdata   => pulse_90deg_s1_readdata,                --                    .readdata
			out_port   => pulse_90deg_external_connection_export  -- external_connection.export
		);

	pulse_t1 : component soc_system_v5_nmr_parameters_delay_t1
		port map (
			clk        => pulse_t1_clk_clk,                    --                 clk.clk
			reset_n    => pulse_t1_reset_reset_n,              --               reset.reset_n
			address    => pulse_t1_s1_address,                 --                  s1.address
			write_n    => pulse_t1_s1_write_n,                 --                    .write_n
			writedata  => pulse_t1_s1_writedata,               --                    .writedata
			chipselect => pulse_t1_s1_chipselect,              --                    .chipselect
			readdata   => pulse_t1_s1_readdata,                --                    .readdata
			out_port   => pulse_t1_external_connection_export  -- external_connection.export
		);

	rx_delay : component soc_system_v5_nmr_parameters_delay_t1
		port map (
			clk        => rx_delay_clk_clk,                    --                 clk.clk
			reset_n    => rx_delay_reset_reset_n,              --               reset.reset_n
			address    => rx_delay_s1_address,                 --                  s1.address
			write_n    => rx_delay_s1_write_n,                 --                    .write_n
			writedata  => rx_delay_s1_writedata,               --                    .writedata
			chipselect => rx_delay_s1_chipselect,              --                    .chipselect
			readdata   => rx_delay_s1_readdata,                --                    .readdata
			out_port   => rx_delay_external_connection_export  -- external_connection.export
		);

	samples_per_echo : component soc_system_v5_nmr_parameters_samples_per_echo
		port map (
			clk        => samples_per_echo_clk_clk,                    --                 clk.clk
			reset_n    => samples_per_echo_reset_reset_n,              --               reset.reset_n
			address    => samples_per_echo_s1_address,                 --                  s1.address
			write_n    => samples_per_echo_s1_write_n,                 --                    .write_n
			writedata  => samples_per_echo_s1_writedata,               --                    .writedata
			chipselect => samples_per_echo_s1_chipselect,              --                    .chipselect
			readdata   => samples_per_echo_s1_readdata,                --                    .readdata
			out_port   => samples_per_echo_external_connection_export  -- external_connection.export
		);

end architecture rtl; -- of soc_system_v5_nmr_parameters
