-- soc_system_v5.vhd

-- Generated using ACDS version 17.1 590

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity soc_system_v5 is
	port (
		adc_fifo_in_data                          : in    std_logic_vector(15 downto 0) := (others => '0'); --                 adc_fifo_in.data
		adc_fifo_in_valid                         : in    std_logic                     := '0';             --                            .valid
		adc_fifo_in_ready                         : out   std_logic;                                        --                            .ready
		adc_val_sub_export                        : out   std_logic_vector(31 downto 0);                    --                 adc_val_sub.export
		alt_vip_itc_0_clocked_video_vid_clk       : in    std_logic                     := '0';             -- alt_vip_itc_0_clocked_video.vid_clk
		alt_vip_itc_0_clocked_video_vid_data      : out   std_logic_vector(31 downto 0);                    --                            .vid_data
		alt_vip_itc_0_clocked_video_underflow     : out   std_logic;                                        --                            .underflow
		alt_vip_itc_0_clocked_video_vid_datavalid : out   std_logic;                                        --                            .vid_datavalid
		alt_vip_itc_0_clocked_video_vid_v_sync    : out   std_logic;                                        --                            .vid_v_sync
		alt_vip_itc_0_clocked_video_vid_h_sync    : out   std_logic;                                        --                            .vid_h_sync
		alt_vip_itc_0_clocked_video_vid_f         : out   std_logic;                                        --                            .vid_f
		alt_vip_itc_0_clocked_video_vid_h         : out   std_logic;                                        --                            .vid_h
		alt_vip_itc_0_clocked_video_vid_v         : out   std_logic;                                        --                            .vid_v
		analyzer_pll_locked_export                : out   std_logic;                                        --         analyzer_pll_locked.export
		analyzer_pll_outclk0_clk                  : out   std_logic;                                        --        analyzer_pll_outclk0.clk
		analyzer_pll_outclk1_clk                  : out   std_logic;                                        --        analyzer_pll_outclk1.clk
		analyzer_pll_outclk2_clk                  : out   std_logic;                                        --        analyzer_pll_outclk2.clk
		analyzer_pll_outclk3_clk                  : out   std_logic;                                        --        analyzer_pll_outclk3.clk
		analyzer_pll_reset_reset                  : in    std_logic                     := '0';             --          analyzer_pll_reset.reset
		aux_cnt_out_export                        : out   std_logic_vector(31 downto 0);                    --                 aux_cnt_out.export
		clk_clk                                   : in    std_logic                     := '0';             --                         clk.clk
		ctrl_in_export                            : in    std_logic_vector(7 downto 0)  := (others => '0'); --                     ctrl_in.export
		ctrl_out_export                           : out   std_logic_vector(31 downto 0);                    --                    ctrl_out.export
		dac_grad_MISO                             : in    std_logic                     := '0';             --                    dac_grad.MISO
		dac_grad_MOSI                             : out   std_logic;                                        --                            .MOSI
		dac_grad_SCLK                             : out   std_logic;                                        --                            .SCLK
		dac_grad_SS_n                             : out   std_logic;                                        --                            .SS_n
		dconv_fifo_in_data                        : in    std_logic_vector(31 downto 0) := (others => '0'); --               dconv_fifo_in.data
		dconv_fifo_in_valid                       : in    std_logic                     := '0';             --                            .valid
		dconv_fifo_in_ready                       : out   std_logic;                                        --                            .ready
		dconv_fifo_q_in_data                      : in    std_logic_vector(31 downto 0) := (others => '0'); --             dconv_fifo_q_in.data
		dconv_fifo_q_in_valid                     : in    std_logic                     := '0';             --                            .valid
		dconv_fifo_q_in_ready                     : out   std_logic;                                        --                            .ready
		dconv_fir_in_data                         : in    std_logic_vector(14 downto 0) := (others => '0'); --                dconv_fir_in.data
		dconv_fir_in_valid                        : in    std_logic                     := '0';             --                            .valid
		dconv_fir_in_error                        : in    std_logic_vector(1 downto 0)  := (others => '0'); --                            .error
		dconv_fir_out_data                        : out   std_logic_vector(31 downto 0);                    --               dconv_fir_out.data
		dconv_fir_out_valid                       : out   std_logic;                                        --                            .valid
		dconv_fir_out_error                       : out   std_logic_vector(1 downto 0);                     --                            .error
		dconv_fir_q_in_data                       : in    std_logic_vector(14 downto 0) := (others => '0'); --              dconv_fir_q_in.data
		dconv_fir_q_in_valid                      : in    std_logic                     := '0';             --                            .valid
		dconv_fir_q_in_error                      : in    std_logic_vector(1 downto 0)  := (others => '0'); --                            .error
		dconv_fir_q_out_data                      : out   std_logic_vector(31 downto 0);                    --             dconv_fir_q_out.data
		dconv_fir_q_out_valid                     : out   std_logic;                                        --                            .valid
		dconv_fir_q_out_error                     : out   std_logic_vector(1 downto 0);                     --                            .error
		delay_nosig_export                        : out   std_logic_vector(31 downto 0);                    --                 delay_nosig.export
		delay_sig_export                          : out   std_logic_vector(31 downto 0);                    --                   delay_sig.export
		delay_t1_export                           : out   std_logic_vector(31 downto 0);                    --                    delay_t1.export
		echoes_per_scan_export                    : out   std_logic_vector(31 downto 0);                    --             echoes_per_scan.export
		fifo_clk_bridge_in_clk                    : in    std_logic                     := '0';             --          fifo_clk_bridge_in.clk
		fifo_rst_reset                            : in    std_logic                     := '0';             --                    fifo_rst.reset
		hps_0_h2f_reset_reset_n                   : out   std_logic;                                        --             hps_0_h2f_reset.reset_n
		hps_0_hps_io_hps_io_emac1_inst_TX_CLK     : out   std_logic;                                        --                hps_0_hps_io.hps_io_emac1_inst_TX_CLK
		hps_0_hps_io_hps_io_emac1_inst_TXD0       : out   std_logic;                                        --                            .hps_io_emac1_inst_TXD0
		hps_0_hps_io_hps_io_emac1_inst_TXD1       : out   std_logic;                                        --                            .hps_io_emac1_inst_TXD1
		hps_0_hps_io_hps_io_emac1_inst_TXD2       : out   std_logic;                                        --                            .hps_io_emac1_inst_TXD2
		hps_0_hps_io_hps_io_emac1_inst_TXD3       : out   std_logic;                                        --                            .hps_io_emac1_inst_TXD3
		hps_0_hps_io_hps_io_emac1_inst_RXD0       : in    std_logic                     := '0';             --                            .hps_io_emac1_inst_RXD0
		hps_0_hps_io_hps_io_emac1_inst_MDIO       : inout std_logic                     := '0';             --                            .hps_io_emac1_inst_MDIO
		hps_0_hps_io_hps_io_emac1_inst_MDC        : out   std_logic;                                        --                            .hps_io_emac1_inst_MDC
		hps_0_hps_io_hps_io_emac1_inst_RX_CTL     : in    std_logic                     := '0';             --                            .hps_io_emac1_inst_RX_CTL
		hps_0_hps_io_hps_io_emac1_inst_TX_CTL     : out   std_logic;                                        --                            .hps_io_emac1_inst_TX_CTL
		hps_0_hps_io_hps_io_emac1_inst_RX_CLK     : in    std_logic                     := '0';             --                            .hps_io_emac1_inst_RX_CLK
		hps_0_hps_io_hps_io_emac1_inst_RXD1       : in    std_logic                     := '0';             --                            .hps_io_emac1_inst_RXD1
		hps_0_hps_io_hps_io_emac1_inst_RXD2       : in    std_logic                     := '0';             --                            .hps_io_emac1_inst_RXD2
		hps_0_hps_io_hps_io_emac1_inst_RXD3       : in    std_logic                     := '0';             --                            .hps_io_emac1_inst_RXD3
		hps_0_hps_io_hps_io_qspi_inst_IO0         : inout std_logic                     := '0';             --                            .hps_io_qspi_inst_IO0
		hps_0_hps_io_hps_io_qspi_inst_IO1         : inout std_logic                     := '0';             --                            .hps_io_qspi_inst_IO1
		hps_0_hps_io_hps_io_qspi_inst_IO2         : inout std_logic                     := '0';             --                            .hps_io_qspi_inst_IO2
		hps_0_hps_io_hps_io_qspi_inst_IO3         : inout std_logic                     := '0';             --                            .hps_io_qspi_inst_IO3
		hps_0_hps_io_hps_io_qspi_inst_SS0         : out   std_logic;                                        --                            .hps_io_qspi_inst_SS0
		hps_0_hps_io_hps_io_qspi_inst_CLK         : out   std_logic;                                        --                            .hps_io_qspi_inst_CLK
		hps_0_hps_io_hps_io_sdio_inst_CMD         : inout std_logic                     := '0';             --                            .hps_io_sdio_inst_CMD
		hps_0_hps_io_hps_io_sdio_inst_D0          : inout std_logic                     := '0';             --                            .hps_io_sdio_inst_D0
		hps_0_hps_io_hps_io_sdio_inst_D1          : inout std_logic                     := '0';             --                            .hps_io_sdio_inst_D1
		hps_0_hps_io_hps_io_sdio_inst_CLK         : out   std_logic;                                        --                            .hps_io_sdio_inst_CLK
		hps_0_hps_io_hps_io_sdio_inst_D2          : inout std_logic                     := '0';             --                            .hps_io_sdio_inst_D2
		hps_0_hps_io_hps_io_sdio_inst_D3          : inout std_logic                     := '0';             --                            .hps_io_sdio_inst_D3
		hps_0_hps_io_hps_io_usb1_inst_D0          : inout std_logic                     := '0';             --                            .hps_io_usb1_inst_D0
		hps_0_hps_io_hps_io_usb1_inst_D1          : inout std_logic                     := '0';             --                            .hps_io_usb1_inst_D1
		hps_0_hps_io_hps_io_usb1_inst_D2          : inout std_logic                     := '0';             --                            .hps_io_usb1_inst_D2
		hps_0_hps_io_hps_io_usb1_inst_D3          : inout std_logic                     := '0';             --                            .hps_io_usb1_inst_D3
		hps_0_hps_io_hps_io_usb1_inst_D4          : inout std_logic                     := '0';             --                            .hps_io_usb1_inst_D4
		hps_0_hps_io_hps_io_usb1_inst_D5          : inout std_logic                     := '0';             --                            .hps_io_usb1_inst_D5
		hps_0_hps_io_hps_io_usb1_inst_D6          : inout std_logic                     := '0';             --                            .hps_io_usb1_inst_D6
		hps_0_hps_io_hps_io_usb1_inst_D7          : inout std_logic                     := '0';             --                            .hps_io_usb1_inst_D7
		hps_0_hps_io_hps_io_usb1_inst_CLK         : in    std_logic                     := '0';             --                            .hps_io_usb1_inst_CLK
		hps_0_hps_io_hps_io_usb1_inst_STP         : out   std_logic;                                        --                            .hps_io_usb1_inst_STP
		hps_0_hps_io_hps_io_usb1_inst_DIR         : in    std_logic                     := '0';             --                            .hps_io_usb1_inst_DIR
		hps_0_hps_io_hps_io_usb1_inst_NXT         : in    std_logic                     := '0';             --                            .hps_io_usb1_inst_NXT
		hps_0_hps_io_hps_io_spim1_inst_CLK        : out   std_logic;                                        --                            .hps_io_spim1_inst_CLK
		hps_0_hps_io_hps_io_spim1_inst_MOSI       : out   std_logic;                                        --                            .hps_io_spim1_inst_MOSI
		hps_0_hps_io_hps_io_spim1_inst_MISO       : in    std_logic                     := '0';             --                            .hps_io_spim1_inst_MISO
		hps_0_hps_io_hps_io_spim1_inst_SS0        : out   std_logic;                                        --                            .hps_io_spim1_inst_SS0
		hps_0_hps_io_hps_io_uart0_inst_RX         : in    std_logic                     := '0';             --                            .hps_io_uart0_inst_RX
		hps_0_hps_io_hps_io_uart0_inst_TX         : out   std_logic;                                        --                            .hps_io_uart0_inst_TX
		hps_0_hps_io_hps_io_i2c0_inst_SDA         : inout std_logic                     := '0';             --                            .hps_io_i2c0_inst_SDA
		hps_0_hps_io_hps_io_i2c0_inst_SCL         : inout std_logic                     := '0';             --                            .hps_io_i2c0_inst_SCL
		hps_0_hps_io_hps_io_i2c1_inst_SDA         : inout std_logic                     := '0';             --                            .hps_io_i2c1_inst_SDA
		hps_0_hps_io_hps_io_i2c1_inst_SCL         : inout std_logic                     := '0';             --                            .hps_io_i2c1_inst_SCL
		hps_0_hps_io_hps_io_gpio_inst_GPIO09      : inout std_logic                     := '0';             --                            .hps_io_gpio_inst_GPIO09
		hps_0_hps_io_hps_io_gpio_inst_GPIO35      : inout std_logic                     := '0';             --                            .hps_io_gpio_inst_GPIO35
		hps_0_hps_io_hps_io_gpio_inst_GPIO40      : inout std_logic                     := '0';             --                            .hps_io_gpio_inst_GPIO40
		hps_0_hps_io_hps_io_gpio_inst_GPIO48      : inout std_logic                     := '0';             --                            .hps_io_gpio_inst_GPIO48
		hps_0_hps_io_hps_io_gpio_inst_GPIO53      : inout std_logic                     := '0';             --                            .hps_io_gpio_inst_GPIO53
		hps_0_hps_io_hps_io_gpio_inst_GPIO54      : inout std_logic                     := '0';             --                            .hps_io_gpio_inst_GPIO54
		hps_0_hps_io_hps_io_gpio_inst_GPIO61      : inout std_logic                     := '0';             --                            .hps_io_gpio_inst_GPIO61
		i2c_ext_sda_in                            : in    std_logic                     := '0';             --                     i2c_ext.sda_in
		i2c_ext_scl_in                            : in    std_logic                     := '0';             --                            .scl_in
		i2c_ext_sda_oe                            : out   std_logic;                                        --                            .sda_oe
		i2c_ext_scl_oe                            : out   std_logic;                                        --                            .scl_oe
		i2c_int_sda_in                            : in    std_logic                     := '0';             --                     i2c_int.sda_in
		i2c_int_scl_in                            : in    std_logic                     := '0';             --                            .scl_in
		i2c_int_sda_oe                            : out   std_logic;                                        --                            .sda_oe
		i2c_int_scl_oe                            : out   std_logic;                                        --                            .scl_oe
		init_delay_export                         : out   std_logic_vector(31 downto 0);                    --                  init_delay.export
		memory_mem_a                              : out   std_logic_vector(14 downto 0);                    --                      memory.mem_a
		memory_mem_ba                             : out   std_logic_vector(2 downto 0);                     --                            .mem_ba
		memory_mem_ck                             : out   std_logic;                                        --                            .mem_ck
		memory_mem_ck_n                           : out   std_logic;                                        --                            .mem_ck_n
		memory_mem_cke                            : out   std_logic;                                        --                            .mem_cke
		memory_mem_cs_n                           : out   std_logic;                                        --                            .mem_cs_n
		memory_mem_ras_n                          : out   std_logic;                                        --                            .mem_ras_n
		memory_mem_cas_n                          : out   std_logic;                                        --                            .mem_cas_n
		memory_mem_we_n                           : out   std_logic;                                        --                            .mem_we_n
		memory_mem_reset_n                        : out   std_logic;                                        --                            .mem_reset_n
		memory_mem_dq                             : inout std_logic_vector(31 downto 0) := (others => '0'); --                            .mem_dq
		memory_mem_dqs                            : inout std_logic_vector(3 downto 0)  := (others => '0'); --                            .mem_dqs
		memory_mem_dqs_n                          : inout std_logic_vector(3 downto 0)  := (others => '0'); --                            .mem_dqs_n
		memory_mem_odt                            : out   std_logic;                                        --                            .mem_odt
		memory_mem_dm                             : out   std_logic_vector(3 downto 0);                     --                            .mem_dm
		memory_oct_rzqin                          : in    std_logic                     := '0';             --                            .oct_rzqin
		nmr_sys_pll_locked_export                 : out   std_logic;                                        --          nmr_sys_pll_locked.export
		nmr_sys_pll_outclk_clk                    : out   std_logic;                                        --          nmr_sys_pll_outclk.clk
		nmr_sys_pll_reset_reset                   : in    std_logic                     := '0';             --           nmr_sys_pll_reset.reset
		pll_vga_clk65_clk                         : out   std_logic;                                        --               pll_vga_clk65.clk
		pll_vga_locked_export                     : out   std_logic;                                        --              pll_vga_locked.export
		pulse_180deg_export                       : out   std_logic_vector(31 downto 0);                    --                pulse_180deg.export
		pulse_90deg_export                        : out   std_logic_vector(31 downto 0);                    --                 pulse_90deg.export
		pulse_t1_export                           : out   std_logic_vector(31 downto 0);                    --                    pulse_t1.export
		reset_reset_n                             : in    std_logic                     := '0';             --                       reset.reset_n
		rx_delay_export                           : out   std_logic_vector(31 downto 0);                    --                    rx_delay.export
		samples_per_echo_export                   : out   std_logic_vector(31 downto 0);                    --            samples_per_echo.export
		sdram_clk_clk                             : out   std_logic;                                        --                   sdram_clk.clk
		sdram_wire_addr                           : out   std_logic_vector(12 downto 0);                    --                  sdram_wire.addr
		sdram_wire_ba                             : out   std_logic_vector(1 downto 0);                     --                            .ba
		sdram_wire_cas_n                          : out   std_logic;                                        --                            .cas_n
		sdram_wire_cke                            : out   std_logic;                                        --                            .cke
		sdram_wire_cs_n                           : out   std_logic;                                        --                            .cs_n
		sdram_wire_dq                             : inout std_logic_vector(15 downto 0) := (others => '0'); --                            .dq
		sdram_wire_dqm                            : out   std_logic_vector(1 downto 0);                     --                            .dqm
		sdram_wire_ras_n                          : out   std_logic;                                        --                            .ras_n
		sdram_wire_we_n                           : out   std_logic;                                        --                            .we_n
		spi_afe_relays_MISO                       : in    std_logic                     := '0';             --              spi_afe_relays.MISO
		spi_afe_relays_MOSI                       : out   std_logic;                                        --                            .MOSI
		spi_afe_relays_SCLK                       : out   std_logic;                                        --                            .SCLK
		spi_afe_relays_SS_n                       : out   std_logic;                                        --                            .SS_n
		spi_mtch_ntwrk_MISO                       : in    std_logic                     := '0';             --              spi_mtch_ntwrk.MISO
		spi_mtch_ntwrk_MOSI                       : out   std_logic;                                        --                            .MOSI
		spi_mtch_ntwrk_SCLK                       : out   std_logic;                                        --                            .SCLK
		spi_mtch_ntwrk_SS_n                       : out   std_logic;                                        --                            .SS_n
		switches_export                           : in    std_logic_vector(9 downto 0)  := (others => '0')  --                    switches.export
	);
end entity soc_system_v5;

architecture rtl of soc_system_v5 is
	component soc_system_v5_adc_fifo_mem is
		port (
			wrclock                         : in  std_logic                     := 'X';             -- clk
			reset_n                         : in  std_logic                     := 'X';             -- reset_n
			avalonst_sink_valid             : in  std_logic                     := 'X';             -- valid
			avalonst_sink_data              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			avalonst_sink_ready             : out std_logic;                                        -- ready
			avalonmm_read_slave_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			avalonmm_read_slave_read        : in  std_logic                     := 'X';             -- read
			avalonmm_read_slave_address     : in  std_logic                     := 'X';             -- address
			avalonmm_read_slave_waitrequest : out std_logic;                                        -- waitrequest
			wrclk_control_slave_address     : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			wrclk_control_slave_read        : in  std_logic                     := 'X';             -- read
			wrclk_control_slave_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			wrclk_control_slave_write       : in  std_logic                     := 'X';             -- write
			wrclk_control_slave_readdata    : out std_logic_vector(31 downto 0)                     -- readdata
		);
	end component soc_system_v5_adc_fifo_mem;

	component soc_system_v5_alt_vip_itc_0 is
		port (
			is_clk        : in  std_logic                     := 'X';             -- clk
			rst           : in  std_logic                     := 'X';             -- reset
			is_data       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			is_valid      : in  std_logic                     := 'X';             -- valid
			is_ready      : out std_logic;                                        -- ready
			is_sop        : in  std_logic                     := 'X';             -- startofpacket
			is_eop        : in  std_logic                     := 'X';             -- endofpacket
			vid_clk       : in  std_logic                     := 'X';             -- export
			vid_data      : out std_logic_vector(31 downto 0);                    -- export
			underflow     : out std_logic;                                        -- export
			vid_datavalid : out std_logic;                                        -- export
			vid_v_sync    : out std_logic;                                        -- export
			vid_h_sync    : out std_logic;                                        -- export
			vid_f         : out std_logic;                                        -- export
			vid_h         : out std_logic;                                        -- export
			vid_v         : out std_logic                                         -- export
		);
	end component soc_system_v5_alt_vip_itc_0;

	component soc_system_v5_alt_vip_vfr_vga is
		port (
			clock                : in  std_logic                      := 'X';             -- clk
			reset                : in  std_logic                      := 'X';             -- reset
			master_clock         : in  std_logic                      := 'X';             -- clk
			master_reset         : in  std_logic                      := 'X';             -- reset
			slave_address        : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- address
			slave_write          : in  std_logic                      := 'X';             -- write
			slave_writedata      : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			slave_read           : in  std_logic                      := 'X';             -- read
			slave_readdata       : out std_logic_vector(31 downto 0);                     -- readdata
			slave_irq            : out std_logic;                                         -- irq
			dout_data            : out std_logic_vector(31 downto 0);                     -- data
			dout_valid           : out std_logic;                                         -- valid
			dout_ready           : in  std_logic                      := 'X';             -- ready
			dout_startofpacket   : out std_logic;                                         -- startofpacket
			dout_endofpacket     : out std_logic;                                         -- endofpacket
			master_address       : out std_logic_vector(31 downto 0);                     -- address
			master_burstcount    : out std_logic_vector(5 downto 0);                      -- burstcount
			master_readdata      : in  std_logic_vector(127 downto 0) := (others => 'X'); -- readdata
			master_read          : out std_logic;                                         -- read
			master_readdatavalid : in  std_logic                      := 'X';             -- readdatavalid
			master_waitrequest   : in  std_logic                      := 'X'              -- waitrequest
		);
	end component soc_system_v5_alt_vip_vfr_vga;

	component soc_system_v5_analyzer_pll is
		port (
			refclk            : in  std_logic                     := 'X';             -- clk
			rst               : in  std_logic                     := 'X';             -- reset
			outclk_0          : out std_logic;                                        -- clk
			outclk_1          : out std_logic;                                        -- clk
			outclk_2          : out std_logic;                                        -- clk
			outclk_3          : out std_logic;                                        -- clk
			locked            : out std_logic;                                        -- export
			reconfig_to_pll   : in  std_logic_vector(63 downto 0) := (others => 'X'); -- reconfig_to_pll
			reconfig_from_pll : out std_logic_vector(63 downto 0)                     -- reconfig_from_pll
		);
	end component soc_system_v5_analyzer_pll;

	component altera_pll_reconfig_top is
		generic (
			device_family       : string  := "";
			ENABLE_MIF          : boolean := false;
			MIF_FILE_NAME       : string  := "";
			ENABLE_BYTEENABLE   : boolean := false;
			BYTEENABLE_WIDTH    : integer := 4;
			RECONFIG_ADDR_WIDTH : integer := 6;
			RECONFIG_DATA_WIDTH : integer := 32;
			reconf_width        : integer := 64;
			WAIT_FOR_LOCK       : boolean := true
		);
		port (
			mgmt_clk          : in  std_logic                     := 'X';             -- clk
			mgmt_reset        : in  std_logic                     := 'X';             -- reset
			mgmt_waitrequest  : out std_logic;                                        -- waitrequest
			mgmt_read         : in  std_logic                     := 'X';             -- read
			mgmt_write        : in  std_logic                     := 'X';             -- write
			mgmt_readdata     : out std_logic_vector(31 downto 0);                    -- readdata
			mgmt_address      : in  std_logic_vector(5 downto 0)  := (others => 'X'); -- address
			mgmt_writedata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			reconfig_to_pll   : out std_logic_vector(63 downto 0);                    -- reconfig_to_pll
			reconfig_from_pll : in  std_logic_vector(63 downto 0) := (others => 'X'); -- reconfig_from_pll
			mgmt_byteenable   : in  std_logic_vector(3 downto 0)  := (others => 'X')  -- byteenable
		);
	end component altera_pll_reconfig_top;

	component soc_system_v5_aux_cnt_out is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(31 downto 0)                     -- export
		);
	end component soc_system_v5_aux_cnt_out;

	component soc_system_v5_ctrl_in is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(7 downto 0)  := (others => 'X')  -- export
		);
	end component soc_system_v5_ctrl_in;

	component soc_system_v5_dac_grad is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			data_from_cpu : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			data_to_cpu   : out std_logic_vector(31 downto 0);                    -- readdata
			mem_addr      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			read_n        : in  std_logic                     := 'X';             -- read_n
			spi_select    : in  std_logic                     := 'X';             -- chipselect
			write_n       : in  std_logic                     := 'X';             -- write_n
			irq           : out std_logic;                                        -- irq
			MISO          : in  std_logic                     := 'X';             -- export
			MOSI          : out std_logic;                                        -- export
			SCLK          : out std_logic;                                        -- export
			SS_n          : out std_logic                                         -- export
		);
	end component soc_system_v5_dac_grad;

	component soc_system_v5_dconv_fifo_mem is
		port (
			wrclock                         : in  std_logic                     := 'X';             -- clk
			reset_n                         : in  std_logic                     := 'X';             -- reset_n
			avalonst_sink_valid             : in  std_logic                     := 'X';             -- valid
			avalonst_sink_data              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			avalonst_sink_ready             : out std_logic;                                        -- ready
			avalonmm_read_slave_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			avalonmm_read_slave_read        : in  std_logic                     := 'X';             -- read
			avalonmm_read_slave_address     : in  std_logic                     := 'X';             -- address
			avalonmm_read_slave_waitrequest : out std_logic;                                        -- waitrequest
			wrclk_control_slave_address     : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			wrclk_control_slave_read        : in  std_logic                     := 'X';             -- read
			wrclk_control_slave_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			wrclk_control_slave_write       : in  std_logic                     := 'X';             -- write
			wrclk_control_slave_readdata    : out std_logic_vector(31 downto 0)                     -- readdata
		);
	end component soc_system_v5_dconv_fifo_mem;

	component soc_system_v5_dconv_fir is
		port (
			clk              : in  std_logic                     := 'X';             -- clk
			reset_n          : in  std_logic                     := 'X';             -- reset_n
			ast_sink_data    : in  std_logic_vector(14 downto 0) := (others => 'X'); -- data
			ast_sink_valid   : in  std_logic                     := 'X';             -- valid
			ast_sink_error   : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- error
			ast_source_data  : out std_logic_vector(31 downto 0);                    -- data
			ast_source_valid : out std_logic;                                        -- valid
			ast_source_error : out std_logic_vector(1 downto 0);                     -- error
			coeff_in_clk     : in  std_logic                     := 'X';             -- clk
			coeff_in_areset  : in  std_logic                     := 'X';             -- reset_n
			coeff_in_address : in  std_logic_vector(5 downto 0)  := (others => 'X'); -- address
			coeff_in_read    : in  std_logic                     := 'X';             -- read
			coeff_out_valid  : out std_logic_vector(0 downto 0);                     -- readdatavalid
			coeff_out_data   : out std_logic_vector(15 downto 0);                    -- readdata
			coeff_in_we      : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- write
			coeff_in_data    : in  std_logic_vector(15 downto 0) := (others => 'X')  -- writedata
		);
	end component soc_system_v5_dconv_fir;

	component soc_system_v5_dma_dconvi is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			system_reset_n     : in  std_logic                     := 'X';             -- reset_n
			dma_ctl_address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			dma_ctl_chipselect : in  std_logic                     := 'X';             -- chipselect
			dma_ctl_readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			dma_ctl_write_n    : in  std_logic                     := 'X';             -- write_n
			dma_ctl_writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dma_ctl_irq        : out std_logic;                                        -- irq
			read_address       : out std_logic_vector(10 downto 0);                    -- address
			read_chipselect    : out std_logic;                                        -- chipselect
			read_read_n        : out std_logic;                                        -- read_n
			read_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			read_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			read_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			write_address      : out std_logic_vector(25 downto 0);                    -- address
			write_chipselect   : out std_logic;                                        -- chipselect
			write_waitrequest  : in  std_logic                     := 'X';             -- waitrequest
			write_write_n      : out std_logic;                                        -- write_n
			write_writedata    : out std_logic_vector(31 downto 0);                    -- writedata
			write_byteenable   : out std_logic_vector(3 downto 0)                      -- byteenable
		);
	end component soc_system_v5_dma_dconvi;

	component soc_system_v5_dma_dconvq is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			system_reset_n     : in  std_logic                     := 'X';             -- reset_n
			dma_ctl_address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			dma_ctl_chipselect : in  std_logic                     := 'X';             -- chipselect
			dma_ctl_readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			dma_ctl_write_n    : in  std_logic                     := 'X';             -- write_n
			dma_ctl_writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dma_ctl_irq        : out std_logic;                                        -- irq
			read_address       : out std_logic_vector(10 downto 0);                    -- address
			read_chipselect    : out std_logic;                                        -- chipselect
			read_read_n        : out std_logic;                                        -- read_n
			read_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			read_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			read_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			write_address      : out std_logic_vector(25 downto 0);                    -- address
			write_chipselect   : out std_logic;                                        -- chipselect
			write_waitrequest  : in  std_logic                     := 'X';             -- waitrequest
			write_write_n      : out std_logic;                                        -- write_n
			write_writedata    : out std_logic_vector(31 downto 0);                    -- writedata
			write_byteenable   : out std_logic_vector(3 downto 0)                      -- byteenable
		);
	end component soc_system_v5_dma_dconvq;

	component soc_system_v5_dma_dummy is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			system_reset_n     : in  std_logic                     := 'X';             -- reset_n
			dma_ctl_address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			dma_ctl_chipselect : in  std_logic                     := 'X';             -- chipselect
			dma_ctl_readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			dma_ctl_write_n    : in  std_logic                     := 'X';             -- write_n
			dma_ctl_writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dma_ctl_irq        : out std_logic;                                        -- irq
			read_address       : out std_logic_vector(26 downto 0);                    -- address
			read_chipselect    : out std_logic;                                        -- chipselect
			read_read_n        : out std_logic;                                        -- read_n
			read_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			read_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			read_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			write_address      : out std_logic_vector(25 downto 0);                    -- address
			write_chipselect   : out std_logic;                                        -- chipselect
			write_waitrequest  : in  std_logic                     := 'X';             -- waitrequest
			write_write_n      : out std_logic;                                        -- write_n
			write_writedata    : out std_logic_vector(31 downto 0);                    -- writedata
			write_byteenable   : out std_logic_vector(3 downto 0)                      -- byteenable
		);
	end component soc_system_v5_dma_dummy;

	component soc_system_v5_dma_fifo is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			system_reset_n     : in  std_logic                     := 'X';             -- reset_n
			dma_ctl_address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			dma_ctl_chipselect : in  std_logic                     := 'X';             -- chipselect
			dma_ctl_readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			dma_ctl_write_n    : in  std_logic                     := 'X';             -- write_n
			dma_ctl_writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dma_ctl_irq        : out std_logic;                                        -- irq
			read_address       : out std_logic_vector(26 downto 0);                    -- address
			read_chipselect    : out std_logic;                                        -- chipselect
			read_read_n        : out std_logic;                                        -- read_n
			read_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			read_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			read_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			write_address      : out std_logic_vector(25 downto 0);                    -- address
			write_chipselect   : out std_logic;                                        -- chipselect
			write_waitrequest  : in  std_logic                     := 'X';             -- waitrequest
			write_write_n      : out std_logic;                                        -- write_n
			write_writedata    : out std_logic_vector(31 downto 0);                    -- writedata
			write_byteenable   : out std_logic_vector(3 downto 0)                      -- byteenable
		);
	end component soc_system_v5_dma_fifo;

	component soc_system_v5_fifo_dummy is
		port (
			wrclock                          : in  std_logic                     := 'X';             -- clk
			reset_n                          : in  std_logic                     := 'X';             -- reset_n
			avalonmm_write_slave_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avalonmm_write_slave_write       : in  std_logic                     := 'X';             -- write
			avalonmm_write_slave_waitrequest : out std_logic;                                        -- waitrequest
			avalonmm_read_slave_readdata     : out std_logic_vector(31 downto 0);                    -- readdata
			avalonmm_read_slave_read         : in  std_logic                     := 'X';             -- read
			avalonmm_read_slave_waitrequest  : out std_logic;                                        -- waitrequest
			wrclk_control_slave_address      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			wrclk_control_slave_read         : in  std_logic                     := 'X';             -- read
			wrclk_control_slave_writedata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			wrclk_control_slave_write        : in  std_logic                     := 'X';             -- write
			wrclk_control_slave_readdata     : out std_logic_vector(31 downto 0)                     -- readdata
		);
	end component soc_system_v5_fifo_dummy;

	component soc_system_v5_fifo_dummy64_in is
		port (
			wrclock                          : in  std_logic                     := 'X';             -- clk
			reset_n                          : in  std_logic                     := 'X';             -- reset_n
			avalonmm_write_slave_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avalonmm_write_slave_write       : in  std_logic                     := 'X';             -- write
			avalonmm_write_slave_address     : in  std_logic                     := 'X';             -- address
			avalonmm_write_slave_waitrequest : out std_logic;                                        -- waitrequest
			avalonst_source_valid            : out std_logic;                                        -- valid
			avalonst_source_data             : out std_logic_vector(31 downto 0);                    -- data
			avalonst_source_ready            : in  std_logic                     := 'X';             -- ready
			wrclk_control_slave_address      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			wrclk_control_slave_read         : in  std_logic                     := 'X';             -- read
			wrclk_control_slave_writedata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			wrclk_control_slave_write        : in  std_logic                     := 'X';             -- write
			wrclk_control_slave_readdata     : out std_logic_vector(31 downto 0)                     -- readdata
		);
	end component soc_system_v5_fifo_dummy64_in;

	component soc_system_v5_fifo_dummy64_out is
		port (
			wrclock                         : in  std_logic                     := 'X';             -- clk
			reset_n                         : in  std_logic                     := 'X';             -- reset_n
			avalonst_sink_valid             : in  std_logic                     := 'X';             -- valid
			avalonst_sink_data              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			avalonst_sink_ready             : out std_logic;                                        -- ready
			avalonmm_read_slave_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			avalonmm_read_slave_read        : in  std_logic                     := 'X';             -- read
			avalonmm_read_slave_address     : in  std_logic                     := 'X';             -- address
			avalonmm_read_slave_waitrequest : out std_logic;                                        -- waitrequest
			wrclk_control_slave_address     : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			wrclk_control_slave_read        : in  std_logic                     := 'X';             -- read
			wrclk_control_slave_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			wrclk_control_slave_write       : in  std_logic                     := 'X';             -- write
			wrclk_control_slave_readdata    : out std_logic_vector(31 downto 0)                     -- readdata
		);
	end component soc_system_v5_fifo_dummy64_out;

	component soc_system_v5_gp_pll is
		port (
			refclk   : in  std_logic := 'X'; -- clk
			rst      : in  std_logic := 'X'; -- reset
			outclk_0 : out std_logic;        -- clk
			outclk_1 : out std_logic;        -- clk
			outclk_2 : out std_logic;        -- clk
			outclk_3 : out std_logic;        -- clk
			locked   : out std_logic         -- export
		);
	end component soc_system_v5_gp_pll;

	component soc_system_v5_hps_0 is
		generic (
			F2S_Width : integer := 2;
			S2F_Width : integer := 2
		);
		port (
			mem_a                    : out   std_logic_vector(14 downto 0);                     -- mem_a
			mem_ba                   : out   std_logic_vector(2 downto 0);                      -- mem_ba
			mem_ck                   : out   std_logic;                                         -- mem_ck
			mem_ck_n                 : out   std_logic;                                         -- mem_ck_n
			mem_cke                  : out   std_logic;                                         -- mem_cke
			mem_cs_n                 : out   std_logic;                                         -- mem_cs_n
			mem_ras_n                : out   std_logic;                                         -- mem_ras_n
			mem_cas_n                : out   std_logic;                                         -- mem_cas_n
			mem_we_n                 : out   std_logic;                                         -- mem_we_n
			mem_reset_n              : out   std_logic;                                         -- mem_reset_n
			mem_dq                   : inout std_logic_vector(31 downto 0)  := (others => 'X'); -- mem_dq
			mem_dqs                  : inout std_logic_vector(3 downto 0)   := (others => 'X'); -- mem_dqs
			mem_dqs_n                : inout std_logic_vector(3 downto 0)   := (others => 'X'); -- mem_dqs_n
			mem_odt                  : out   std_logic;                                         -- mem_odt
			mem_dm                   : out   std_logic_vector(3 downto 0);                      -- mem_dm
			oct_rzqin                : in    std_logic                      := 'X';             -- oct_rzqin
			hps_io_emac1_inst_TX_CLK : out   std_logic;                                         -- hps_io_emac1_inst_TX_CLK
			hps_io_emac1_inst_TXD0   : out   std_logic;                                         -- hps_io_emac1_inst_TXD0
			hps_io_emac1_inst_TXD1   : out   std_logic;                                         -- hps_io_emac1_inst_TXD1
			hps_io_emac1_inst_TXD2   : out   std_logic;                                         -- hps_io_emac1_inst_TXD2
			hps_io_emac1_inst_TXD3   : out   std_logic;                                         -- hps_io_emac1_inst_TXD3
			hps_io_emac1_inst_RXD0   : in    std_logic                      := 'X';             -- hps_io_emac1_inst_RXD0
			hps_io_emac1_inst_MDIO   : inout std_logic                      := 'X';             -- hps_io_emac1_inst_MDIO
			hps_io_emac1_inst_MDC    : out   std_logic;                                         -- hps_io_emac1_inst_MDC
			hps_io_emac1_inst_RX_CTL : in    std_logic                      := 'X';             -- hps_io_emac1_inst_RX_CTL
			hps_io_emac1_inst_TX_CTL : out   std_logic;                                         -- hps_io_emac1_inst_TX_CTL
			hps_io_emac1_inst_RX_CLK : in    std_logic                      := 'X';             -- hps_io_emac1_inst_RX_CLK
			hps_io_emac1_inst_RXD1   : in    std_logic                      := 'X';             -- hps_io_emac1_inst_RXD1
			hps_io_emac1_inst_RXD2   : in    std_logic                      := 'X';             -- hps_io_emac1_inst_RXD2
			hps_io_emac1_inst_RXD3   : in    std_logic                      := 'X';             -- hps_io_emac1_inst_RXD3
			hps_io_qspi_inst_IO0     : inout std_logic                      := 'X';             -- hps_io_qspi_inst_IO0
			hps_io_qspi_inst_IO1     : inout std_logic                      := 'X';             -- hps_io_qspi_inst_IO1
			hps_io_qspi_inst_IO2     : inout std_logic                      := 'X';             -- hps_io_qspi_inst_IO2
			hps_io_qspi_inst_IO3     : inout std_logic                      := 'X';             -- hps_io_qspi_inst_IO3
			hps_io_qspi_inst_SS0     : out   std_logic;                                         -- hps_io_qspi_inst_SS0
			hps_io_qspi_inst_CLK     : out   std_logic;                                         -- hps_io_qspi_inst_CLK
			hps_io_sdio_inst_CMD     : inout std_logic                      := 'X';             -- hps_io_sdio_inst_CMD
			hps_io_sdio_inst_D0      : inout std_logic                      := 'X';             -- hps_io_sdio_inst_D0
			hps_io_sdio_inst_D1      : inout std_logic                      := 'X';             -- hps_io_sdio_inst_D1
			hps_io_sdio_inst_CLK     : out   std_logic;                                         -- hps_io_sdio_inst_CLK
			hps_io_sdio_inst_D2      : inout std_logic                      := 'X';             -- hps_io_sdio_inst_D2
			hps_io_sdio_inst_D3      : inout std_logic                      := 'X';             -- hps_io_sdio_inst_D3
			hps_io_usb1_inst_D0      : inout std_logic                      := 'X';             -- hps_io_usb1_inst_D0
			hps_io_usb1_inst_D1      : inout std_logic                      := 'X';             -- hps_io_usb1_inst_D1
			hps_io_usb1_inst_D2      : inout std_logic                      := 'X';             -- hps_io_usb1_inst_D2
			hps_io_usb1_inst_D3      : inout std_logic                      := 'X';             -- hps_io_usb1_inst_D3
			hps_io_usb1_inst_D4      : inout std_logic                      := 'X';             -- hps_io_usb1_inst_D4
			hps_io_usb1_inst_D5      : inout std_logic                      := 'X';             -- hps_io_usb1_inst_D5
			hps_io_usb1_inst_D6      : inout std_logic                      := 'X';             -- hps_io_usb1_inst_D6
			hps_io_usb1_inst_D7      : inout std_logic                      := 'X';             -- hps_io_usb1_inst_D7
			hps_io_usb1_inst_CLK     : in    std_logic                      := 'X';             -- hps_io_usb1_inst_CLK
			hps_io_usb1_inst_STP     : out   std_logic;                                         -- hps_io_usb1_inst_STP
			hps_io_usb1_inst_DIR     : in    std_logic                      := 'X';             -- hps_io_usb1_inst_DIR
			hps_io_usb1_inst_NXT     : in    std_logic                      := 'X';             -- hps_io_usb1_inst_NXT
			hps_io_spim1_inst_CLK    : out   std_logic;                                         -- hps_io_spim1_inst_CLK
			hps_io_spim1_inst_MOSI   : out   std_logic;                                         -- hps_io_spim1_inst_MOSI
			hps_io_spim1_inst_MISO   : in    std_logic                      := 'X';             -- hps_io_spim1_inst_MISO
			hps_io_spim1_inst_SS0    : out   std_logic;                                         -- hps_io_spim1_inst_SS0
			hps_io_uart0_inst_RX     : in    std_logic                      := 'X';             -- hps_io_uart0_inst_RX
			hps_io_uart0_inst_TX     : out   std_logic;                                         -- hps_io_uart0_inst_TX
			hps_io_i2c0_inst_SDA     : inout std_logic                      := 'X';             -- hps_io_i2c0_inst_SDA
			hps_io_i2c0_inst_SCL     : inout std_logic                      := 'X';             -- hps_io_i2c0_inst_SCL
			hps_io_i2c1_inst_SDA     : inout std_logic                      := 'X';             -- hps_io_i2c1_inst_SDA
			hps_io_i2c1_inst_SCL     : inout std_logic                      := 'X';             -- hps_io_i2c1_inst_SCL
			hps_io_gpio_inst_GPIO09  : inout std_logic                      := 'X';             -- hps_io_gpio_inst_GPIO09
			hps_io_gpio_inst_GPIO35  : inout std_logic                      := 'X';             -- hps_io_gpio_inst_GPIO35
			hps_io_gpio_inst_GPIO40  : inout std_logic                      := 'X';             -- hps_io_gpio_inst_GPIO40
			hps_io_gpio_inst_GPIO48  : inout std_logic                      := 'X';             -- hps_io_gpio_inst_GPIO48
			hps_io_gpio_inst_GPIO53  : inout std_logic                      := 'X';             -- hps_io_gpio_inst_GPIO53
			hps_io_gpio_inst_GPIO54  : inout std_logic                      := 'X';             -- hps_io_gpio_inst_GPIO54
			hps_io_gpio_inst_GPIO61  : inout std_logic                      := 'X';             -- hps_io_gpio_inst_GPIO61
			h2f_rst_n                : out   std_logic;                                         -- reset_n
			h2f_axi_clk              : in    std_logic                      := 'X';             -- clk
			h2f_AWID                 : out   std_logic_vector(11 downto 0);                     -- awid
			h2f_AWADDR               : out   std_logic_vector(29 downto 0);                     -- awaddr
			h2f_AWLEN                : out   std_logic_vector(3 downto 0);                      -- awlen
			h2f_AWSIZE               : out   std_logic_vector(2 downto 0);                      -- awsize
			h2f_AWBURST              : out   std_logic_vector(1 downto 0);                      -- awburst
			h2f_AWLOCK               : out   std_logic_vector(1 downto 0);                      -- awlock
			h2f_AWCACHE              : out   std_logic_vector(3 downto 0);                      -- awcache
			h2f_AWPROT               : out   std_logic_vector(2 downto 0);                      -- awprot
			h2f_AWVALID              : out   std_logic;                                         -- awvalid
			h2f_AWREADY              : in    std_logic                      := 'X';             -- awready
			h2f_WID                  : out   std_logic_vector(11 downto 0);                     -- wid
			h2f_WDATA                : out   std_logic_vector(127 downto 0);                    -- wdata
			h2f_WSTRB                : out   std_logic_vector(15 downto 0);                     -- wstrb
			h2f_WLAST                : out   std_logic;                                         -- wlast
			h2f_WVALID               : out   std_logic;                                         -- wvalid
			h2f_WREADY               : in    std_logic                      := 'X';             -- wready
			h2f_BID                  : in    std_logic_vector(11 downto 0)  := (others => 'X'); -- bid
			h2f_BRESP                : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- bresp
			h2f_BVALID               : in    std_logic                      := 'X';             -- bvalid
			h2f_BREADY               : out   std_logic;                                         -- bready
			h2f_ARID                 : out   std_logic_vector(11 downto 0);                     -- arid
			h2f_ARADDR               : out   std_logic_vector(29 downto 0);                     -- araddr
			h2f_ARLEN                : out   std_logic_vector(3 downto 0);                      -- arlen
			h2f_ARSIZE               : out   std_logic_vector(2 downto 0);                      -- arsize
			h2f_ARBURST              : out   std_logic_vector(1 downto 0);                      -- arburst
			h2f_ARLOCK               : out   std_logic_vector(1 downto 0);                      -- arlock
			h2f_ARCACHE              : out   std_logic_vector(3 downto 0);                      -- arcache
			h2f_ARPROT               : out   std_logic_vector(2 downto 0);                      -- arprot
			h2f_ARVALID              : out   std_logic;                                         -- arvalid
			h2f_ARREADY              : in    std_logic                      := 'X';             -- arready
			h2f_RID                  : in    std_logic_vector(11 downto 0)  := (others => 'X'); -- rid
			h2f_RDATA                : in    std_logic_vector(127 downto 0) := (others => 'X'); -- rdata
			h2f_RRESP                : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- rresp
			h2f_RLAST                : in    std_logic                      := 'X';             -- rlast
			h2f_RVALID               : in    std_logic                      := 'X';             -- rvalid
			h2f_RREADY               : out   std_logic;                                         -- rready
			f2h_axi_clk              : in    std_logic                      := 'X';             -- clk
			f2h_AWID                 : in    std_logic_vector(7 downto 0)   := (others => 'X'); -- awid
			f2h_AWADDR               : in    std_logic_vector(31 downto 0)  := (others => 'X'); -- awaddr
			f2h_AWLEN                : in    std_logic_vector(3 downto 0)   := (others => 'X'); -- awlen
			f2h_AWSIZE               : in    std_logic_vector(2 downto 0)   := (others => 'X'); -- awsize
			f2h_AWBURST              : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- awburst
			f2h_AWLOCK               : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- awlock
			f2h_AWCACHE              : in    std_logic_vector(3 downto 0)   := (others => 'X'); -- awcache
			f2h_AWPROT               : in    std_logic_vector(2 downto 0)   := (others => 'X'); -- awprot
			f2h_AWVALID              : in    std_logic                      := 'X';             -- awvalid
			f2h_AWREADY              : out   std_logic;                                         -- awready
			f2h_AWUSER               : in    std_logic_vector(4 downto 0)   := (others => 'X'); -- awuser
			f2h_WID                  : in    std_logic_vector(7 downto 0)   := (others => 'X'); -- wid
			f2h_WDATA                : in    std_logic_vector(127 downto 0) := (others => 'X'); -- wdata
			f2h_WSTRB                : in    std_logic_vector(15 downto 0)  := (others => 'X'); -- wstrb
			f2h_WLAST                : in    std_logic                      := 'X';             -- wlast
			f2h_WVALID               : in    std_logic                      := 'X';             -- wvalid
			f2h_WREADY               : out   std_logic;                                         -- wready
			f2h_BID                  : out   std_logic_vector(7 downto 0);                      -- bid
			f2h_BRESP                : out   std_logic_vector(1 downto 0);                      -- bresp
			f2h_BVALID               : out   std_logic;                                         -- bvalid
			f2h_BREADY               : in    std_logic                      := 'X';             -- bready
			f2h_ARID                 : in    std_logic_vector(7 downto 0)   := (others => 'X'); -- arid
			f2h_ARADDR               : in    std_logic_vector(31 downto 0)  := (others => 'X'); -- araddr
			f2h_ARLEN                : in    std_logic_vector(3 downto 0)   := (others => 'X'); -- arlen
			f2h_ARSIZE               : in    std_logic_vector(2 downto 0)   := (others => 'X'); -- arsize
			f2h_ARBURST              : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- arburst
			f2h_ARLOCK               : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- arlock
			f2h_ARCACHE              : in    std_logic_vector(3 downto 0)   := (others => 'X'); -- arcache
			f2h_ARPROT               : in    std_logic_vector(2 downto 0)   := (others => 'X'); -- arprot
			f2h_ARVALID              : in    std_logic                      := 'X';             -- arvalid
			f2h_ARREADY              : out   std_logic;                                         -- arready
			f2h_ARUSER               : in    std_logic_vector(4 downto 0)   := (others => 'X'); -- aruser
			f2h_RID                  : out   std_logic_vector(7 downto 0);                      -- rid
			f2h_RDATA                : out   std_logic_vector(127 downto 0);                    -- rdata
			f2h_RRESP                : out   std_logic_vector(1 downto 0);                      -- rresp
			f2h_RLAST                : out   std_logic;                                         -- rlast
			f2h_RVALID               : out   std_logic;                                         -- rvalid
			f2h_RREADY               : in    std_logic                      := 'X';             -- rready
			h2f_lw_axi_clk           : in    std_logic                      := 'X';             -- clk
			h2f_lw_AWID              : out   std_logic_vector(11 downto 0);                     -- awid
			h2f_lw_AWADDR            : out   std_logic_vector(20 downto 0);                     -- awaddr
			h2f_lw_AWLEN             : out   std_logic_vector(3 downto 0);                      -- awlen
			h2f_lw_AWSIZE            : out   std_logic_vector(2 downto 0);                      -- awsize
			h2f_lw_AWBURST           : out   std_logic_vector(1 downto 0);                      -- awburst
			h2f_lw_AWLOCK            : out   std_logic_vector(1 downto 0);                      -- awlock
			h2f_lw_AWCACHE           : out   std_logic_vector(3 downto 0);                      -- awcache
			h2f_lw_AWPROT            : out   std_logic_vector(2 downto 0);                      -- awprot
			h2f_lw_AWVALID           : out   std_logic;                                         -- awvalid
			h2f_lw_AWREADY           : in    std_logic                      := 'X';             -- awready
			h2f_lw_WID               : out   std_logic_vector(11 downto 0);                     -- wid
			h2f_lw_WDATA             : out   std_logic_vector(31 downto 0);                     -- wdata
			h2f_lw_WSTRB             : out   std_logic_vector(3 downto 0);                      -- wstrb
			h2f_lw_WLAST             : out   std_logic;                                         -- wlast
			h2f_lw_WVALID            : out   std_logic;                                         -- wvalid
			h2f_lw_WREADY            : in    std_logic                      := 'X';             -- wready
			h2f_lw_BID               : in    std_logic_vector(11 downto 0)  := (others => 'X'); -- bid
			h2f_lw_BRESP             : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- bresp
			h2f_lw_BVALID            : in    std_logic                      := 'X';             -- bvalid
			h2f_lw_BREADY            : out   std_logic;                                         -- bready
			h2f_lw_ARID              : out   std_logic_vector(11 downto 0);                     -- arid
			h2f_lw_ARADDR            : out   std_logic_vector(20 downto 0);                     -- araddr
			h2f_lw_ARLEN             : out   std_logic_vector(3 downto 0);                      -- arlen
			h2f_lw_ARSIZE            : out   std_logic_vector(2 downto 0);                      -- arsize
			h2f_lw_ARBURST           : out   std_logic_vector(1 downto 0);                      -- arburst
			h2f_lw_ARLOCK            : out   std_logic_vector(1 downto 0);                      -- arlock
			h2f_lw_ARCACHE           : out   std_logic_vector(3 downto 0);                      -- arcache
			h2f_lw_ARPROT            : out   std_logic_vector(2 downto 0);                      -- arprot
			h2f_lw_ARVALID           : out   std_logic;                                         -- arvalid
			h2f_lw_ARREADY           : in    std_logic                      := 'X';             -- arready
			h2f_lw_RID               : in    std_logic_vector(11 downto 0)  := (others => 'X'); -- rid
			h2f_lw_RDATA             : in    std_logic_vector(31 downto 0)  := (others => 'X'); -- rdata
			h2f_lw_RRESP             : in    std_logic_vector(1 downto 0)   := (others => 'X'); -- rresp
			h2f_lw_RLAST             : in    std_logic                      := 'X';             -- rlast
			h2f_lw_RVALID            : in    std_logic                      := 'X';             -- rvalid
			h2f_lw_RREADY            : out   std_logic;                                         -- rready
			f2h_irq_p0               : in    std_logic_vector(31 downto 0)  := (others => 'X'); -- irq
			f2h_irq_p1               : in    std_logic_vector(31 downto 0)  := (others => 'X')  -- irq
		);
	end component soc_system_v5_hps_0;

	component altera_avalon_i2c is
		generic (
			USE_AV_ST       : integer := 0;
			FIFO_DEPTH      : integer := 4;
			FIFO_DEPTH_LOG2 : integer := 2
		);
		port (
			clk       : in  std_logic                     := 'X';             -- clk
			rst_n     : in  std_logic                     := 'X';             -- reset_n
			intr      : out std_logic;                                        -- irq
			addr      : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- address
			read      : in  std_logic                     := 'X';             -- read
			write     : in  std_logic                     := 'X';             -- write
			writedata : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata  : out std_logic_vector(31 downto 0);                    -- readdata
			sda_in    : in  std_logic                     := 'X';             -- sda_in
			scl_in    : in  std_logic                     := 'X';             -- scl_in
			sda_oe    : out std_logic;                                        -- sda_oe
			scl_oe    : out std_logic;                                        -- scl_oe
			src_data  : out std_logic_vector(7 downto 0);                     -- data
			src_valid : out std_logic;                                        -- valid
			src_ready : in  std_logic                     := 'X';             -- ready
			snk_data  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- data
			snk_valid : in  std_logic                     := 'X';             -- valid
			snk_ready : out std_logic                                         -- ready
		);
	end component altera_avalon_i2c;

	component soc_system_v5_jtag_uart is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component soc_system_v5_jtag_uart;

	component soc_system_v5_master_non_sec is
		generic (
			USE_PLI     : integer := 0;
			PLI_PORT    : integer := 50000;
			FIFO_DEPTHS : integer := 2
		);
		port (
			clk_clk              : in  std_logic                     := 'X';             -- clk
			clk_reset_reset      : in  std_logic                     := 'X';             -- reset
			master_address       : out std_logic_vector(31 downto 0);                    -- address
			master_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			master_read          : out std_logic;                                        -- read
			master_write         : out std_logic;                                        -- write
			master_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			master_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			master_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			master_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			master_reset_reset   : out std_logic                                         -- reset
		);
	end component soc_system_v5_master_non_sec;

	component soc_system_v5_nmr_parameters is
		port (
			adc_val_sub_clk_clk                         : in  std_logic                     := 'X';             -- clk
			adc_val_sub_external_connection_export      : out std_logic_vector(31 downto 0);                    -- export
			adc_val_sub_reset_reset_n                   : in  std_logic                     := 'X';             -- reset_n
			adc_val_sub_s1_address                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			adc_val_sub_s1_write_n                      : in  std_logic                     := 'X';             -- write_n
			adc_val_sub_s1_writedata                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			adc_val_sub_s1_chipselect                   : in  std_logic                     := 'X';             -- chipselect
			adc_val_sub_s1_readdata                     : out std_logic_vector(31 downto 0);                    -- readdata
			delay_nosig_clk_clk                         : in  std_logic                     := 'X';             -- clk
			delay_nosig_external_connection_export      : out std_logic_vector(31 downto 0);                    -- export
			delay_nosig_reset_reset_n                   : in  std_logic                     := 'X';             -- reset_n
			delay_nosig_s1_address                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			delay_nosig_s1_write_n                      : in  std_logic                     := 'X';             -- write_n
			delay_nosig_s1_writedata                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			delay_nosig_s1_chipselect                   : in  std_logic                     := 'X';             -- chipselect
			delay_nosig_s1_readdata                     : out std_logic_vector(31 downto 0);                    -- readdata
			delay_sig_clk_clk                           : in  std_logic                     := 'X';             -- clk
			delay_sig_external_connection_export        : out std_logic_vector(31 downto 0);                    -- export
			delay_sig_reset_reset_n                     : in  std_logic                     := 'X';             -- reset_n
			delay_sig_s1_address                        : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			delay_sig_s1_write_n                        : in  std_logic                     := 'X';             -- write_n
			delay_sig_s1_writedata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			delay_sig_s1_chipselect                     : in  std_logic                     := 'X';             -- chipselect
			delay_sig_s1_readdata                       : out std_logic_vector(31 downto 0);                    -- readdata
			delay_t1_clk_clk                            : in  std_logic                     := 'X';             -- clk
			delay_t1_external_connection_export         : out std_logic_vector(31 downto 0);                    -- export
			delay_t1_reset_reset_n                      : in  std_logic                     := 'X';             -- reset_n
			delay_t1_s1_address                         : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			delay_t1_s1_write_n                         : in  std_logic                     := 'X';             -- write_n
			delay_t1_s1_writedata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			delay_t1_s1_chipselect                      : in  std_logic                     := 'X';             -- chipselect
			delay_t1_s1_readdata                        : out std_logic_vector(31 downto 0);                    -- readdata
			echoes_per_scan_clk_clk                     : in  std_logic                     := 'X';             -- clk
			echoes_per_scan_external_connection_export  : out std_logic_vector(31 downto 0);                    -- export
			echoes_per_scan_reset_reset_n               : in  std_logic                     := 'X';             -- reset_n
			echoes_per_scan_s1_address                  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			echoes_per_scan_s1_write_n                  : in  std_logic                     := 'X';             -- write_n
			echoes_per_scan_s1_writedata                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			echoes_per_scan_s1_chipselect               : in  std_logic                     := 'X';             -- chipselect
			echoes_per_scan_s1_readdata                 : out std_logic_vector(31 downto 0);                    -- readdata
			init_delay_clk_clk                          : in  std_logic                     := 'X';             -- clk
			init_delay_external_connection_export       : out std_logic_vector(31 downto 0);                    -- export
			init_delay_reset_reset_n                    : in  std_logic                     := 'X';             -- reset_n
			init_delay_s1_address                       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			init_delay_s1_write_n                       : in  std_logic                     := 'X';             -- write_n
			init_delay_s1_writedata                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			init_delay_s1_chipselect                    : in  std_logic                     := 'X';             -- chipselect
			init_delay_s1_readdata                      : out std_logic_vector(31 downto 0);                    -- readdata
			pulse_180deg_clk_clk                        : in  std_logic                     := 'X';             -- clk
			pulse_180deg_external_connection_export     : out std_logic_vector(31 downto 0);                    -- export
			pulse_180deg_reset_reset_n                  : in  std_logic                     := 'X';             -- reset_n
			pulse_180deg_s1_address                     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			pulse_180deg_s1_write_n                     : in  std_logic                     := 'X';             -- write_n
			pulse_180deg_s1_writedata                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			pulse_180deg_s1_chipselect                  : in  std_logic                     := 'X';             -- chipselect
			pulse_180deg_s1_readdata                    : out std_logic_vector(31 downto 0);                    -- readdata
			pulse_90deg_clk_clk                         : in  std_logic                     := 'X';             -- clk
			pulse_90deg_external_connection_export      : out std_logic_vector(31 downto 0);                    -- export
			pulse_90deg_reset_reset_n                   : in  std_logic                     := 'X';             -- reset_n
			pulse_90deg_s1_address                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			pulse_90deg_s1_write_n                      : in  std_logic                     := 'X';             -- write_n
			pulse_90deg_s1_writedata                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			pulse_90deg_s1_chipselect                   : in  std_logic                     := 'X';             -- chipselect
			pulse_90deg_s1_readdata                     : out std_logic_vector(31 downto 0);                    -- readdata
			pulse_t1_clk_clk                            : in  std_logic                     := 'X';             -- clk
			pulse_t1_external_connection_export         : out std_logic_vector(31 downto 0);                    -- export
			pulse_t1_reset_reset_n                      : in  std_logic                     := 'X';             -- reset_n
			pulse_t1_s1_address                         : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			pulse_t1_s1_write_n                         : in  std_logic                     := 'X';             -- write_n
			pulse_t1_s1_writedata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			pulse_t1_s1_chipselect                      : in  std_logic                     := 'X';             -- chipselect
			pulse_t1_s1_readdata                        : out std_logic_vector(31 downto 0);                    -- readdata
			rx_delay_clk_clk                            : in  std_logic                     := 'X';             -- clk
			rx_delay_external_connection_export         : out std_logic_vector(31 downto 0);                    -- export
			rx_delay_reset_reset_n                      : in  std_logic                     := 'X';             -- reset_n
			rx_delay_s1_address                         : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			rx_delay_s1_write_n                         : in  std_logic                     := 'X';             -- write_n
			rx_delay_s1_writedata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			rx_delay_s1_chipselect                      : in  std_logic                     := 'X';             -- chipselect
			rx_delay_s1_readdata                        : out std_logic_vector(31 downto 0);                    -- readdata
			samples_per_echo_clk_clk                    : in  std_logic                     := 'X';             -- clk
			samples_per_echo_external_connection_export : out std_logic_vector(31 downto 0);                    -- export
			samples_per_echo_reset_reset_n              : in  std_logic                     := 'X';             -- reset_n
			samples_per_echo_s1_address                 : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			samples_per_echo_s1_write_n                 : in  std_logic                     := 'X';             -- write_n
			samples_per_echo_s1_writedata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			samples_per_echo_s1_chipselect              : in  std_logic                     := 'X';             -- chipselect
			samples_per_echo_s1_readdata                : out std_logic_vector(31 downto 0)                     -- readdata
		);
	end component soc_system_v5_nmr_parameters;

	component soc_system_v5_nmr_sys_pll is
		port (
			refclk            : in  std_logic                     := 'X';             -- clk
			rst               : in  std_logic                     := 'X';             -- reset
			outclk_0          : out std_logic;                                        -- clk
			locked            : out std_logic;                                        -- export
			reconfig_to_pll   : in  std_logic_vector(63 downto 0) := (others => 'X'); -- reconfig_to_pll
			reconfig_from_pll : out std_logic_vector(63 downto 0)                     -- reconfig_from_pll
		);
	end component soc_system_v5_nmr_sys_pll;

	component soc_system_v5_sdram is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(24 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(12 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component soc_system_v5_sdram;

	component soc_system_v5_spi_afe_relays is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			data_from_cpu : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			data_to_cpu   : out std_logic_vector(31 downto 0);                    -- readdata
			mem_addr      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			read_n        : in  std_logic                     := 'X';             -- read_n
			spi_select    : in  std_logic                     := 'X';             -- chipselect
			write_n       : in  std_logic                     := 'X';             -- write_n
			irq           : out std_logic;                                        -- irq
			MISO          : in  std_logic                     := 'X';             -- export
			MOSI          : out std_logic;                                        -- export
			SCLK          : out std_logic;                                        -- export
			SS_n          : out std_logic                                         -- export
		);
	end component soc_system_v5_spi_afe_relays;

	component soc_system_v5_switches is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(9 downto 0)  := (others => 'X')  -- export
		);
	end component soc_system_v5_switches;

	component soc_system_v5_sysid_qsys is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component soc_system_v5_sysid_qsys;

	component soc_system_v5_mm_interconnect_0 is
		port (
			hps_0_f2h_axi_slave_awid                                         : out std_logic_vector(7 downto 0);                      -- awid
			hps_0_f2h_axi_slave_awaddr                                       : out std_logic_vector(31 downto 0);                     -- awaddr
			hps_0_f2h_axi_slave_awlen                                        : out std_logic_vector(3 downto 0);                      -- awlen
			hps_0_f2h_axi_slave_awsize                                       : out std_logic_vector(2 downto 0);                      -- awsize
			hps_0_f2h_axi_slave_awburst                                      : out std_logic_vector(1 downto 0);                      -- awburst
			hps_0_f2h_axi_slave_awlock                                       : out std_logic_vector(1 downto 0);                      -- awlock
			hps_0_f2h_axi_slave_awcache                                      : out std_logic_vector(3 downto 0);                      -- awcache
			hps_0_f2h_axi_slave_awprot                                       : out std_logic_vector(2 downto 0);                      -- awprot
			hps_0_f2h_axi_slave_awuser                                       : out std_logic_vector(4 downto 0);                      -- awuser
			hps_0_f2h_axi_slave_awvalid                                      : out std_logic;                                         -- awvalid
			hps_0_f2h_axi_slave_awready                                      : in  std_logic                      := 'X';             -- awready
			hps_0_f2h_axi_slave_wid                                          : out std_logic_vector(7 downto 0);                      -- wid
			hps_0_f2h_axi_slave_wdata                                        : out std_logic_vector(127 downto 0);                    -- wdata
			hps_0_f2h_axi_slave_wstrb                                        : out std_logic_vector(15 downto 0);                     -- wstrb
			hps_0_f2h_axi_slave_wlast                                        : out std_logic;                                         -- wlast
			hps_0_f2h_axi_slave_wvalid                                       : out std_logic;                                         -- wvalid
			hps_0_f2h_axi_slave_wready                                       : in  std_logic                      := 'X';             -- wready
			hps_0_f2h_axi_slave_bid                                          : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- bid
			hps_0_f2h_axi_slave_bresp                                        : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- bresp
			hps_0_f2h_axi_slave_bvalid                                       : in  std_logic                      := 'X';             -- bvalid
			hps_0_f2h_axi_slave_bready                                       : out std_logic;                                         -- bready
			hps_0_f2h_axi_slave_arid                                         : out std_logic_vector(7 downto 0);                      -- arid
			hps_0_f2h_axi_slave_araddr                                       : out std_logic_vector(31 downto 0);                     -- araddr
			hps_0_f2h_axi_slave_arlen                                        : out std_logic_vector(3 downto 0);                      -- arlen
			hps_0_f2h_axi_slave_arsize                                       : out std_logic_vector(2 downto 0);                      -- arsize
			hps_0_f2h_axi_slave_arburst                                      : out std_logic_vector(1 downto 0);                      -- arburst
			hps_0_f2h_axi_slave_arlock                                       : out std_logic_vector(1 downto 0);                      -- arlock
			hps_0_f2h_axi_slave_arcache                                      : out std_logic_vector(3 downto 0);                      -- arcache
			hps_0_f2h_axi_slave_arprot                                       : out std_logic_vector(2 downto 0);                      -- arprot
			hps_0_f2h_axi_slave_aruser                                       : out std_logic_vector(4 downto 0);                      -- aruser
			hps_0_f2h_axi_slave_arvalid                                      : out std_logic;                                         -- arvalid
			hps_0_f2h_axi_slave_arready                                      : in  std_logic                      := 'X';             -- arready
			hps_0_f2h_axi_slave_rid                                          : in  std_logic_vector(7 downto 0)   := (others => 'X'); -- rid
			hps_0_f2h_axi_slave_rdata                                        : in  std_logic_vector(127 downto 0) := (others => 'X'); -- rdata
			hps_0_f2h_axi_slave_rresp                                        : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- rresp
			hps_0_f2h_axi_slave_rlast                                        : in  std_logic                      := 'X';             -- rlast
			hps_0_f2h_axi_slave_rvalid                                       : in  std_logic                      := 'X';             -- rvalid
			hps_0_f2h_axi_slave_rready                                       : out std_logic;                                         -- rready
			clk_0_clk_clk                                                    : in  std_logic                      := 'X';             -- clk
			alt_vip_vfr_vga_clock_master_reset_reset_bridge_in_reset_reset   : in  std_logic                      := 'X';             -- reset
			hps_0_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset_reset : in  std_logic                      := 'X';             -- reset
			master_secure_clk_reset_reset_bridge_in_reset_reset              : in  std_logic                      := 'X';             -- reset
			alt_vip_vfr_vga_avalon_master_address                            : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- address
			alt_vip_vfr_vga_avalon_master_waitrequest                        : out std_logic;                                         -- waitrequest
			alt_vip_vfr_vga_avalon_master_burstcount                         : in  std_logic_vector(5 downto 0)   := (others => 'X'); -- burstcount
			alt_vip_vfr_vga_avalon_master_read                               : in  std_logic                      := 'X';             -- read
			alt_vip_vfr_vga_avalon_master_readdata                           : out std_logic_vector(127 downto 0);                    -- readdata
			alt_vip_vfr_vga_avalon_master_readdatavalid                      : out std_logic;                                         -- readdatavalid
			master_secure_master_address                                     : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- address
			master_secure_master_waitrequest                                 : out std_logic;                                         -- waitrequest
			master_secure_master_byteenable                                  : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			master_secure_master_read                                        : in  std_logic                      := 'X';             -- read
			master_secure_master_readdata                                    : out std_logic_vector(31 downto 0);                     -- readdata
			master_secure_master_readdatavalid                               : out std_logic;                                         -- readdatavalid
			master_secure_master_write                                       : in  std_logic                      := 'X';             -- write
			master_secure_master_writedata                                   : in  std_logic_vector(31 downto 0)  := (others => 'X')  -- writedata
		);
	end component soc_system_v5_mm_interconnect_0;

	component soc_system_v5_mm_interconnect_1 is
		port (
			hps_0_h2f_axi_master_awid                                        : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- awid
			hps_0_h2f_axi_master_awaddr                                      : in  std_logic_vector(29 downto 0)  := (others => 'X'); -- awaddr
			hps_0_h2f_axi_master_awlen                                       : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- awlen
			hps_0_h2f_axi_master_awsize                                      : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- awsize
			hps_0_h2f_axi_master_awburst                                     : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- awburst
			hps_0_h2f_axi_master_awlock                                      : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- awlock
			hps_0_h2f_axi_master_awcache                                     : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- awcache
			hps_0_h2f_axi_master_awprot                                      : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- awprot
			hps_0_h2f_axi_master_awvalid                                     : in  std_logic                      := 'X';             -- awvalid
			hps_0_h2f_axi_master_awready                                     : out std_logic;                                         -- awready
			hps_0_h2f_axi_master_wid                                         : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- wid
			hps_0_h2f_axi_master_wdata                                       : in  std_logic_vector(127 downto 0) := (others => 'X'); -- wdata
			hps_0_h2f_axi_master_wstrb                                       : in  std_logic_vector(15 downto 0)  := (others => 'X'); -- wstrb
			hps_0_h2f_axi_master_wlast                                       : in  std_logic                      := 'X';             -- wlast
			hps_0_h2f_axi_master_wvalid                                      : in  std_logic                      := 'X';             -- wvalid
			hps_0_h2f_axi_master_wready                                      : out std_logic;                                         -- wready
			hps_0_h2f_axi_master_bid                                         : out std_logic_vector(11 downto 0);                     -- bid
			hps_0_h2f_axi_master_bresp                                       : out std_logic_vector(1 downto 0);                      -- bresp
			hps_0_h2f_axi_master_bvalid                                      : out std_logic;                                         -- bvalid
			hps_0_h2f_axi_master_bready                                      : in  std_logic                      := 'X';             -- bready
			hps_0_h2f_axi_master_arid                                        : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- arid
			hps_0_h2f_axi_master_araddr                                      : in  std_logic_vector(29 downto 0)  := (others => 'X'); -- araddr
			hps_0_h2f_axi_master_arlen                                       : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- arlen
			hps_0_h2f_axi_master_arsize                                      : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- arsize
			hps_0_h2f_axi_master_arburst                                     : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- arburst
			hps_0_h2f_axi_master_arlock                                      : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- arlock
			hps_0_h2f_axi_master_arcache                                     : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- arcache
			hps_0_h2f_axi_master_arprot                                      : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- arprot
			hps_0_h2f_axi_master_arvalid                                     : in  std_logic                      := 'X';             -- arvalid
			hps_0_h2f_axi_master_arready                                     : out std_logic;                                         -- arready
			hps_0_h2f_axi_master_rid                                         : out std_logic_vector(11 downto 0);                     -- rid
			hps_0_h2f_axi_master_rdata                                       : out std_logic_vector(127 downto 0);                    -- rdata
			hps_0_h2f_axi_master_rresp                                       : out std_logic_vector(1 downto 0);                      -- rresp
			hps_0_h2f_axi_master_rlast                                       : out std_logic;                                         -- rlast
			hps_0_h2f_axi_master_rvalid                                      : out std_logic;                                         -- rvalid
			hps_0_h2f_axi_master_rready                                      : in  std_logic                      := 'X';             -- rready
			hps_0_h2f_lw_axi_master_awid                                     : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- awid
			hps_0_h2f_lw_axi_master_awaddr                                   : in  std_logic_vector(20 downto 0)  := (others => 'X'); -- awaddr
			hps_0_h2f_lw_axi_master_awlen                                    : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- awlen
			hps_0_h2f_lw_axi_master_awsize                                   : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- awsize
			hps_0_h2f_lw_axi_master_awburst                                  : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- awburst
			hps_0_h2f_lw_axi_master_awlock                                   : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- awlock
			hps_0_h2f_lw_axi_master_awcache                                  : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- awcache
			hps_0_h2f_lw_axi_master_awprot                                   : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- awprot
			hps_0_h2f_lw_axi_master_awvalid                                  : in  std_logic                      := 'X';             -- awvalid
			hps_0_h2f_lw_axi_master_awready                                  : out std_logic;                                         -- awready
			hps_0_h2f_lw_axi_master_wid                                      : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- wid
			hps_0_h2f_lw_axi_master_wdata                                    : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- wdata
			hps_0_h2f_lw_axi_master_wstrb                                    : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- wstrb
			hps_0_h2f_lw_axi_master_wlast                                    : in  std_logic                      := 'X';             -- wlast
			hps_0_h2f_lw_axi_master_wvalid                                   : in  std_logic                      := 'X';             -- wvalid
			hps_0_h2f_lw_axi_master_wready                                   : out std_logic;                                         -- wready
			hps_0_h2f_lw_axi_master_bid                                      : out std_logic_vector(11 downto 0);                     -- bid
			hps_0_h2f_lw_axi_master_bresp                                    : out std_logic_vector(1 downto 0);                      -- bresp
			hps_0_h2f_lw_axi_master_bvalid                                   : out std_logic;                                         -- bvalid
			hps_0_h2f_lw_axi_master_bready                                   : in  std_logic                      := 'X';             -- bready
			hps_0_h2f_lw_axi_master_arid                                     : in  std_logic_vector(11 downto 0)  := (others => 'X'); -- arid
			hps_0_h2f_lw_axi_master_araddr                                   : in  std_logic_vector(20 downto 0)  := (others => 'X'); -- araddr
			hps_0_h2f_lw_axi_master_arlen                                    : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- arlen
			hps_0_h2f_lw_axi_master_arsize                                   : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- arsize
			hps_0_h2f_lw_axi_master_arburst                                  : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- arburst
			hps_0_h2f_lw_axi_master_arlock                                   : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- arlock
			hps_0_h2f_lw_axi_master_arcache                                  : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- arcache
			hps_0_h2f_lw_axi_master_arprot                                   : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- arprot
			hps_0_h2f_lw_axi_master_arvalid                                  : in  std_logic                      := 'X';             -- arvalid
			hps_0_h2f_lw_axi_master_arready                                  : out std_logic;                                         -- arready
			hps_0_h2f_lw_axi_master_rid                                      : out std_logic_vector(11 downto 0);                     -- rid
			hps_0_h2f_lw_axi_master_rdata                                    : out std_logic_vector(31 downto 0);                     -- rdata
			hps_0_h2f_lw_axi_master_rresp                                    : out std_logic_vector(1 downto 0);                      -- rresp
			hps_0_h2f_lw_axi_master_rlast                                    : out std_logic;                                         -- rlast
			hps_0_h2f_lw_axi_master_rvalid                                   : out std_logic;                                         -- rvalid
			hps_0_h2f_lw_axi_master_rready                                   : in  std_logic                      := 'X';             -- rready
			clk_0_clk_clk                                                    : in  std_logic                      := 'X';             -- clk
			gp_pll_outclk0_clk                                               : in  std_logic                      := 'X';             -- clk
			adc_fifo_mem_reset_in_reset_bridge_in_reset_reset                : in  std_logic                      := 'X';             -- reset
			alt_vip_vfr_vga_clock_reset_reset_reset_bridge_in_reset_reset    : in  std_logic                      := 'X';             -- reset
			dma_fifo_reset_reset_bridge_in_reset_reset                       : in  std_logic                      := 'X';             -- reset
			hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset : in  std_logic                      := 'X';             -- reset
			master_non_sec_clk_reset_reset_bridge_in_reset_reset             : in  std_logic                      := 'X';             -- reset
			dma_dconvi_read_master_address                                   : in  std_logic_vector(10 downto 0)  := (others => 'X'); -- address
			dma_dconvi_read_master_waitrequest                               : out std_logic;                                         -- waitrequest
			dma_dconvi_read_master_chipselect                                : in  std_logic                      := 'X';             -- chipselect
			dma_dconvi_read_master_read                                      : in  std_logic                      := 'X';             -- read
			dma_dconvi_read_master_readdata                                  : out std_logic_vector(31 downto 0);                     -- readdata
			dma_dconvi_read_master_readdatavalid                             : out std_logic;                                         -- readdatavalid
			dma_dconvi_write_master_address                                  : in  std_logic_vector(25 downto 0)  := (others => 'X'); -- address
			dma_dconvi_write_master_waitrequest                              : out std_logic;                                         -- waitrequest
			dma_dconvi_write_master_byteenable                               : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			dma_dconvi_write_master_chipselect                               : in  std_logic                      := 'X';             -- chipselect
			dma_dconvi_write_master_write                                    : in  std_logic                      := 'X';             -- write
			dma_dconvi_write_master_writedata                                : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			dma_dconvq_read_master_address                                   : in  std_logic_vector(10 downto 0)  := (others => 'X'); -- address
			dma_dconvq_read_master_waitrequest                               : out std_logic;                                         -- waitrequest
			dma_dconvq_read_master_chipselect                                : in  std_logic                      := 'X';             -- chipselect
			dma_dconvq_read_master_read                                      : in  std_logic                      := 'X';             -- read
			dma_dconvq_read_master_readdata                                  : out std_logic_vector(31 downto 0);                     -- readdata
			dma_dconvq_read_master_readdatavalid                             : out std_logic;                                         -- readdatavalid
			dma_dconvq_write_master_address                                  : in  std_logic_vector(25 downto 0)  := (others => 'X'); -- address
			dma_dconvq_write_master_waitrequest                              : out std_logic;                                         -- waitrequest
			dma_dconvq_write_master_byteenable                               : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			dma_dconvq_write_master_chipselect                               : in  std_logic                      := 'X';             -- chipselect
			dma_dconvq_write_master_write                                    : in  std_logic                      := 'X';             -- write
			dma_dconvq_write_master_writedata                                : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			dma_dummy_read_master_address                                    : in  std_logic_vector(26 downto 0)  := (others => 'X'); -- address
			dma_dummy_read_master_waitrequest                                : out std_logic;                                         -- waitrequest
			dma_dummy_read_master_chipselect                                 : in  std_logic                      := 'X';             -- chipselect
			dma_dummy_read_master_read                                       : in  std_logic                      := 'X';             -- read
			dma_dummy_read_master_readdata                                   : out std_logic_vector(31 downto 0);                     -- readdata
			dma_dummy_read_master_readdatavalid                              : out std_logic;                                         -- readdatavalid
			dma_dummy_write_master_address                                   : in  std_logic_vector(25 downto 0)  := (others => 'X'); -- address
			dma_dummy_write_master_waitrequest                               : out std_logic;                                         -- waitrequest
			dma_dummy_write_master_byteenable                                : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			dma_dummy_write_master_chipselect                                : in  std_logic                      := 'X';             -- chipselect
			dma_dummy_write_master_write                                     : in  std_logic                      := 'X';             -- write
			dma_dummy_write_master_writedata                                 : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			dma_fifo_read_master_address                                     : in  std_logic_vector(26 downto 0)  := (others => 'X'); -- address
			dma_fifo_read_master_waitrequest                                 : out std_logic;                                         -- waitrequest
			dma_fifo_read_master_chipselect                                  : in  std_logic                      := 'X';             -- chipselect
			dma_fifo_read_master_read                                        : in  std_logic                      := 'X';             -- read
			dma_fifo_read_master_readdata                                    : out std_logic_vector(31 downto 0);                     -- readdata
			dma_fifo_read_master_readdatavalid                               : out std_logic;                                         -- readdatavalid
			dma_fifo_write_master_address                                    : in  std_logic_vector(25 downto 0)  := (others => 'X'); -- address
			dma_fifo_write_master_waitrequest                                : out std_logic;                                         -- waitrequest
			dma_fifo_write_master_byteenable                                 : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			dma_fifo_write_master_chipselect                                 : in  std_logic                      := 'X';             -- chipselect
			dma_fifo_write_master_write                                      : in  std_logic                      := 'X';             -- write
			dma_fifo_write_master_writedata                                  : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			master_non_sec_master_address                                    : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- address
			master_non_sec_master_waitrequest                                : out std_logic;                                         -- waitrequest
			master_non_sec_master_byteenable                                 : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			master_non_sec_master_read                                       : in  std_logic                      := 'X';             -- read
			master_non_sec_master_readdata                                   : out std_logic_vector(31 downto 0);                     -- readdata
			master_non_sec_master_readdatavalid                              : out std_logic;                                         -- readdatavalid
			master_non_sec_master_write                                      : in  std_logic                      := 'X';             -- write
			master_non_sec_master_writedata                                  : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			adc_fifo_mem_in_csr_address                                      : out std_logic_vector(2 downto 0);                      -- address
			adc_fifo_mem_in_csr_write                                        : out std_logic;                                         -- write
			adc_fifo_mem_in_csr_read                                         : out std_logic;                                         -- read
			adc_fifo_mem_in_csr_readdata                                     : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			adc_fifo_mem_in_csr_writedata                                    : out std_logic_vector(31 downto 0);                     -- writedata
			adc_fifo_mem_out_address                                         : out std_logic_vector(0 downto 0);                      -- address
			adc_fifo_mem_out_read                                            : out std_logic;                                         -- read
			adc_fifo_mem_out_readdata                                        : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			adc_fifo_mem_out_waitrequest                                     : in  std_logic                      := 'X';             -- waitrequest
			alt_vip_vfr_vga_avalon_slave_address                             : out std_logic_vector(4 downto 0);                      -- address
			alt_vip_vfr_vga_avalon_slave_write                               : out std_logic;                                         -- write
			alt_vip_vfr_vga_avalon_slave_read                                : out std_logic;                                         -- read
			alt_vip_vfr_vga_avalon_slave_readdata                            : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			alt_vip_vfr_vga_avalon_slave_writedata                           : out std_logic_vector(31 downto 0);                     -- writedata
			analyzer_pll_reconfig_mgmt_avalon_slave_address                  : out std_logic_vector(5 downto 0);                      -- address
			analyzer_pll_reconfig_mgmt_avalon_slave_write                    : out std_logic;                                         -- write
			analyzer_pll_reconfig_mgmt_avalon_slave_read                     : out std_logic;                                         -- read
			analyzer_pll_reconfig_mgmt_avalon_slave_readdata                 : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			analyzer_pll_reconfig_mgmt_avalon_slave_writedata                : out std_logic_vector(31 downto 0);                     -- writedata
			analyzer_pll_reconfig_mgmt_avalon_slave_waitrequest              : in  std_logic                      := 'X';             -- waitrequest
			aux_cnt_out_s1_address                                           : out std_logic_vector(1 downto 0);                      -- address
			aux_cnt_out_s1_write                                             : out std_logic;                                         -- write
			aux_cnt_out_s1_readdata                                          : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			aux_cnt_out_s1_writedata                                         : out std_logic_vector(31 downto 0);                     -- writedata
			aux_cnt_out_s1_chipselect                                        : out std_logic;                                         -- chipselect
			ctrl_in_s1_address                                               : out std_logic_vector(1 downto 0);                      -- address
			ctrl_in_s1_readdata                                              : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			ctrl_out_s1_address                                              : out std_logic_vector(1 downto 0);                      -- address
			ctrl_out_s1_write                                                : out std_logic;                                         -- write
			ctrl_out_s1_readdata                                             : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			ctrl_out_s1_writedata                                            : out std_logic_vector(31 downto 0);                     -- writedata
			ctrl_out_s1_chipselect                                           : out std_logic;                                         -- chipselect
			dac_grad_spi_control_port_address                                : out std_logic_vector(2 downto 0);                      -- address
			dac_grad_spi_control_port_write                                  : out std_logic;                                         -- write
			dac_grad_spi_control_port_read                                   : out std_logic;                                         -- read
			dac_grad_spi_control_port_readdata                               : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			dac_grad_spi_control_port_writedata                              : out std_logic_vector(31 downto 0);                     -- writedata
			dac_grad_spi_control_port_chipselect                             : out std_logic;                                         -- chipselect
			dconv_fifo_mem_in_csr_address                                    : out std_logic_vector(2 downto 0);                      -- address
			dconv_fifo_mem_in_csr_write                                      : out std_logic;                                         -- write
			dconv_fifo_mem_in_csr_read                                       : out std_logic;                                         -- read
			dconv_fifo_mem_in_csr_readdata                                   : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			dconv_fifo_mem_in_csr_writedata                                  : out std_logic_vector(31 downto 0);                     -- writedata
			dconv_fifo_mem_out_address                                       : out std_logic_vector(0 downto 0);                      -- address
			dconv_fifo_mem_out_read                                          : out std_logic;                                         -- read
			dconv_fifo_mem_out_readdata                                      : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			dconv_fifo_mem_out_waitrequest                                   : in  std_logic                      := 'X';             -- waitrequest
			dconv_fifo_mem_q_in_csr_address                                  : out std_logic_vector(2 downto 0);                      -- address
			dconv_fifo_mem_q_in_csr_write                                    : out std_logic;                                         -- write
			dconv_fifo_mem_q_in_csr_read                                     : out std_logic;                                         -- read
			dconv_fifo_mem_q_in_csr_readdata                                 : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			dconv_fifo_mem_q_in_csr_writedata                                : out std_logic_vector(31 downto 0);                     -- writedata
			dconv_fifo_mem_q_out_address                                     : out std_logic_vector(0 downto 0);                      -- address
			dconv_fifo_mem_q_out_read                                        : out std_logic;                                         -- read
			dconv_fifo_mem_q_out_readdata                                    : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			dconv_fifo_mem_q_out_waitrequest                                 : in  std_logic                      := 'X';             -- waitrequest
			dconv_fir_avalon_mm_slave_address                                : out std_logic_vector(5 downto 0);                      -- address
			dconv_fir_avalon_mm_slave_write                                  : out std_logic;                                         -- write
			dconv_fir_avalon_mm_slave_read                                   : out std_logic;                                         -- read
			dconv_fir_avalon_mm_slave_readdata                               : in  std_logic_vector(15 downto 0)  := (others => 'X'); -- readdata
			dconv_fir_avalon_mm_slave_writedata                              : out std_logic_vector(15 downto 0);                     -- writedata
			dconv_fir_avalon_mm_slave_readdatavalid                          : in  std_logic                      := 'X';             -- readdatavalid
			dconv_fir_q_avalon_mm_slave_address                              : out std_logic_vector(5 downto 0);                      -- address
			dconv_fir_q_avalon_mm_slave_write                                : out std_logic;                                         -- write
			dconv_fir_q_avalon_mm_slave_read                                 : out std_logic;                                         -- read
			dconv_fir_q_avalon_mm_slave_readdata                             : in  std_logic_vector(15 downto 0)  := (others => 'X'); -- readdata
			dconv_fir_q_avalon_mm_slave_writedata                            : out std_logic_vector(15 downto 0);                     -- writedata
			dconv_fir_q_avalon_mm_slave_readdatavalid                        : in  std_logic                      := 'X';             -- readdatavalid
			dma_dconvi_control_port_slave_address                            : out std_logic_vector(2 downto 0);                      -- address
			dma_dconvi_control_port_slave_write                              : out std_logic;                                         -- write
			dma_dconvi_control_port_slave_readdata                           : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			dma_dconvi_control_port_slave_writedata                          : out std_logic_vector(31 downto 0);                     -- writedata
			dma_dconvi_control_port_slave_chipselect                         : out std_logic;                                         -- chipselect
			dma_dconvq_control_port_slave_address                            : out std_logic_vector(2 downto 0);                      -- address
			dma_dconvq_control_port_slave_write                              : out std_logic;                                         -- write
			dma_dconvq_control_port_slave_readdata                           : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			dma_dconvq_control_port_slave_writedata                          : out std_logic_vector(31 downto 0);                     -- writedata
			dma_dconvq_control_port_slave_chipselect                         : out std_logic;                                         -- chipselect
			dma_dummy_control_port_slave_address                             : out std_logic_vector(2 downto 0);                      -- address
			dma_dummy_control_port_slave_write                               : out std_logic;                                         -- write
			dma_dummy_control_port_slave_readdata                            : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			dma_dummy_control_port_slave_writedata                           : out std_logic_vector(31 downto 0);                     -- writedata
			dma_dummy_control_port_slave_chipselect                          : out std_logic;                                         -- chipselect
			dma_fifo_control_port_slave_address                              : out std_logic_vector(2 downto 0);                      -- address
			dma_fifo_control_port_slave_write                                : out std_logic;                                         -- write
			dma_fifo_control_port_slave_readdata                             : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			dma_fifo_control_port_slave_writedata                            : out std_logic_vector(31 downto 0);                     -- writedata
			dma_fifo_control_port_slave_chipselect                           : out std_logic;                                         -- chipselect
			fifo_dummy_in_write                                              : out std_logic;                                         -- write
			fifo_dummy_in_writedata                                          : out std_logic_vector(31 downto 0);                     -- writedata
			fifo_dummy_in_waitrequest                                        : in  std_logic                      := 'X';             -- waitrequest
			fifo_dummy_in_csr_address                                        : out std_logic_vector(2 downto 0);                      -- address
			fifo_dummy_in_csr_write                                          : out std_logic;                                         -- write
			fifo_dummy_in_csr_read                                           : out std_logic;                                         -- read
			fifo_dummy_in_csr_readdata                                       : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			fifo_dummy_in_csr_writedata                                      : out std_logic_vector(31 downto 0);                     -- writedata
			fifo_dummy_out_read                                              : out std_logic;                                         -- read
			fifo_dummy_out_readdata                                          : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			fifo_dummy_out_waitrequest                                       : in  std_logic                      := 'X';             -- waitrequest
			fifo_dummy64_in_in_address                                       : out std_logic_vector(0 downto 0);                      -- address
			fifo_dummy64_in_in_write                                         : out std_logic;                                         -- write
			fifo_dummy64_in_in_writedata                                     : out std_logic_vector(31 downto 0);                     -- writedata
			fifo_dummy64_in_in_waitrequest                                   : in  std_logic                      := 'X';             -- waitrequest
			fifo_dummy64_in_in_csr_address                                   : out std_logic_vector(2 downto 0);                      -- address
			fifo_dummy64_in_in_csr_write                                     : out std_logic;                                         -- write
			fifo_dummy64_in_in_csr_read                                      : out std_logic;                                         -- read
			fifo_dummy64_in_in_csr_readdata                                  : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			fifo_dummy64_in_in_csr_writedata                                 : out std_logic_vector(31 downto 0);                     -- writedata
			fifo_dummy64_out_in_csr_address                                  : out std_logic_vector(2 downto 0);                      -- address
			fifo_dummy64_out_in_csr_write                                    : out std_logic;                                         -- write
			fifo_dummy64_out_in_csr_read                                     : out std_logic;                                         -- read
			fifo_dummy64_out_in_csr_readdata                                 : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			fifo_dummy64_out_in_csr_writedata                                : out std_logic_vector(31 downto 0);                     -- writedata
			fifo_dummy64_out_out_address                                     : out std_logic_vector(0 downto 0);                      -- address
			fifo_dummy64_out_out_read                                        : out std_logic;                                         -- read
			fifo_dummy64_out_out_readdata                                    : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			fifo_dummy64_out_out_waitrequest                                 : in  std_logic                      := 'X';             -- waitrequest
			i2c_ext_csr_address                                              : out std_logic_vector(3 downto 0);                      -- address
			i2c_ext_csr_write                                                : out std_logic;                                         -- write
			i2c_ext_csr_read                                                 : out std_logic;                                         -- read
			i2c_ext_csr_readdata                                             : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			i2c_ext_csr_writedata                                            : out std_logic_vector(31 downto 0);                     -- writedata
			i2c_int_csr_address                                              : out std_logic_vector(3 downto 0);                      -- address
			i2c_int_csr_write                                                : out std_logic;                                         -- write
			i2c_int_csr_read                                                 : out std_logic;                                         -- read
			i2c_int_csr_readdata                                             : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			i2c_int_csr_writedata                                            : out std_logic_vector(31 downto 0);                     -- writedata
			jtag_uart_avalon_jtag_slave_address                              : out std_logic_vector(0 downto 0);                      -- address
			jtag_uart_avalon_jtag_slave_write                                : out std_logic;                                         -- write
			jtag_uart_avalon_jtag_slave_read                                 : out std_logic;                                         -- read
			jtag_uart_avalon_jtag_slave_readdata                             : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			jtag_uart_avalon_jtag_slave_writedata                            : out std_logic_vector(31 downto 0);                     -- writedata
			jtag_uart_avalon_jtag_slave_waitrequest                          : in  std_logic                      := 'X';             -- waitrequest
			jtag_uart_avalon_jtag_slave_chipselect                           : out std_logic;                                         -- chipselect
			nmr_parameters_adc_val_sub_s1_address                            : out std_logic_vector(1 downto 0);                      -- address
			nmr_parameters_adc_val_sub_s1_write                              : out std_logic;                                         -- write
			nmr_parameters_adc_val_sub_s1_readdata                           : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			nmr_parameters_adc_val_sub_s1_writedata                          : out std_logic_vector(31 downto 0);                     -- writedata
			nmr_parameters_adc_val_sub_s1_chipselect                         : out std_logic;                                         -- chipselect
			nmr_parameters_delay_nosig_s1_address                            : out std_logic_vector(1 downto 0);                      -- address
			nmr_parameters_delay_nosig_s1_write                              : out std_logic;                                         -- write
			nmr_parameters_delay_nosig_s1_readdata                           : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			nmr_parameters_delay_nosig_s1_writedata                          : out std_logic_vector(31 downto 0);                     -- writedata
			nmr_parameters_delay_nosig_s1_chipselect                         : out std_logic;                                         -- chipselect
			nmr_parameters_delay_sig_s1_address                              : out std_logic_vector(1 downto 0);                      -- address
			nmr_parameters_delay_sig_s1_write                                : out std_logic;                                         -- write
			nmr_parameters_delay_sig_s1_readdata                             : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			nmr_parameters_delay_sig_s1_writedata                            : out std_logic_vector(31 downto 0);                     -- writedata
			nmr_parameters_delay_sig_s1_chipselect                           : out std_logic;                                         -- chipselect
			nmr_parameters_delay_t1_s1_address                               : out std_logic_vector(1 downto 0);                      -- address
			nmr_parameters_delay_t1_s1_write                                 : out std_logic;                                         -- write
			nmr_parameters_delay_t1_s1_readdata                              : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			nmr_parameters_delay_t1_s1_writedata                             : out std_logic_vector(31 downto 0);                     -- writedata
			nmr_parameters_delay_t1_s1_chipselect                            : out std_logic;                                         -- chipselect
			nmr_parameters_echoes_per_scan_s1_address                        : out std_logic_vector(1 downto 0);                      -- address
			nmr_parameters_echoes_per_scan_s1_write                          : out std_logic;                                         -- write
			nmr_parameters_echoes_per_scan_s1_readdata                       : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			nmr_parameters_echoes_per_scan_s1_writedata                      : out std_logic_vector(31 downto 0);                     -- writedata
			nmr_parameters_echoes_per_scan_s1_chipselect                     : out std_logic;                                         -- chipselect
			nmr_parameters_init_delay_s1_address                             : out std_logic_vector(1 downto 0);                      -- address
			nmr_parameters_init_delay_s1_write                               : out std_logic;                                         -- write
			nmr_parameters_init_delay_s1_readdata                            : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			nmr_parameters_init_delay_s1_writedata                           : out std_logic_vector(31 downto 0);                     -- writedata
			nmr_parameters_init_delay_s1_chipselect                          : out std_logic;                                         -- chipselect
			nmr_parameters_pulse_180deg_s1_address                           : out std_logic_vector(1 downto 0);                      -- address
			nmr_parameters_pulse_180deg_s1_write                             : out std_logic;                                         -- write
			nmr_parameters_pulse_180deg_s1_readdata                          : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			nmr_parameters_pulse_180deg_s1_writedata                         : out std_logic_vector(31 downto 0);                     -- writedata
			nmr_parameters_pulse_180deg_s1_chipselect                        : out std_logic;                                         -- chipselect
			nmr_parameters_pulse_90deg_s1_address                            : out std_logic_vector(1 downto 0);                      -- address
			nmr_parameters_pulse_90deg_s1_write                              : out std_logic;                                         -- write
			nmr_parameters_pulse_90deg_s1_readdata                           : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			nmr_parameters_pulse_90deg_s1_writedata                          : out std_logic_vector(31 downto 0);                     -- writedata
			nmr_parameters_pulse_90deg_s1_chipselect                         : out std_logic;                                         -- chipselect
			nmr_parameters_pulse_t1_s1_address                               : out std_logic_vector(1 downto 0);                      -- address
			nmr_parameters_pulse_t1_s1_write                                 : out std_logic;                                         -- write
			nmr_parameters_pulse_t1_s1_readdata                              : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			nmr_parameters_pulse_t1_s1_writedata                             : out std_logic_vector(31 downto 0);                     -- writedata
			nmr_parameters_pulse_t1_s1_chipselect                            : out std_logic;                                         -- chipselect
			nmr_parameters_rx_delay_s1_address                               : out std_logic_vector(1 downto 0);                      -- address
			nmr_parameters_rx_delay_s1_write                                 : out std_logic;                                         -- write
			nmr_parameters_rx_delay_s1_readdata                              : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			nmr_parameters_rx_delay_s1_writedata                             : out std_logic_vector(31 downto 0);                     -- writedata
			nmr_parameters_rx_delay_s1_chipselect                            : out std_logic;                                         -- chipselect
			nmr_parameters_samples_per_echo_s1_address                       : out std_logic_vector(1 downto 0);                      -- address
			nmr_parameters_samples_per_echo_s1_write                         : out std_logic;                                         -- write
			nmr_parameters_samples_per_echo_s1_readdata                      : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			nmr_parameters_samples_per_echo_s1_writedata                     : out std_logic_vector(31 downto 0);                     -- writedata
			nmr_parameters_samples_per_echo_s1_chipselect                    : out std_logic;                                         -- chipselect
			nmr_sys_pll_reconfig_mgmt_avalon_slave_address                   : out std_logic_vector(5 downto 0);                      -- address
			nmr_sys_pll_reconfig_mgmt_avalon_slave_write                     : out std_logic;                                         -- write
			nmr_sys_pll_reconfig_mgmt_avalon_slave_read                      : out std_logic;                                         -- read
			nmr_sys_pll_reconfig_mgmt_avalon_slave_readdata                  : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			nmr_sys_pll_reconfig_mgmt_avalon_slave_writedata                 : out std_logic_vector(31 downto 0);                     -- writedata
			nmr_sys_pll_reconfig_mgmt_avalon_slave_waitrequest               : in  std_logic                      := 'X';             -- waitrequest
			sdram_s1_address                                                 : out std_logic_vector(24 downto 0);                     -- address
			sdram_s1_write                                                   : out std_logic;                                         -- write
			sdram_s1_read                                                    : out std_logic;                                         -- read
			sdram_s1_readdata                                                : in  std_logic_vector(15 downto 0)  := (others => 'X'); -- readdata
			sdram_s1_writedata                                               : out std_logic_vector(15 downto 0);                     -- writedata
			sdram_s1_byteenable                                              : out std_logic_vector(1 downto 0);                      -- byteenable
			sdram_s1_readdatavalid                                           : in  std_logic                      := 'X';             -- readdatavalid
			sdram_s1_waitrequest                                             : in  std_logic                      := 'X';             -- waitrequest
			sdram_s1_chipselect                                              : out std_logic;                                         -- chipselect
			spi_afe_relays_spi_control_port_address                          : out std_logic_vector(2 downto 0);                      -- address
			spi_afe_relays_spi_control_port_write                            : out std_logic;                                         -- write
			spi_afe_relays_spi_control_port_read                             : out std_logic;                                         -- read
			spi_afe_relays_spi_control_port_readdata                         : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			spi_afe_relays_spi_control_port_writedata                        : out std_logic_vector(31 downto 0);                     -- writedata
			spi_afe_relays_spi_control_port_chipselect                       : out std_logic;                                         -- chipselect
			spi_mtch_ntwrk_spi_control_port_address                          : out std_logic_vector(2 downto 0);                      -- address
			spi_mtch_ntwrk_spi_control_port_write                            : out std_logic;                                         -- write
			spi_mtch_ntwrk_spi_control_port_read                             : out std_logic;                                         -- read
			spi_mtch_ntwrk_spi_control_port_readdata                         : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			spi_mtch_ntwrk_spi_control_port_writedata                        : out std_logic_vector(31 downto 0);                     -- writedata
			spi_mtch_ntwrk_spi_control_port_chipselect                       : out std_logic;                                         -- chipselect
			switches_s1_address                                              : out std_logic_vector(1 downto 0);                      -- address
			switches_s1_readdata                                             : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			sysid_qsys_control_slave_address                                 : out std_logic_vector(0 downto 0);                      -- address
			sysid_qsys_control_slave_readdata                                : in  std_logic_vector(31 downto 0)  := (others => 'X')  -- readdata
		);
	end component soc_system_v5_mm_interconnect_1;

	component soc_system_v5_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component soc_system_v5_irq_mapper;

	component soc_system_v5_irq_mapper_001 is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			receiver3_irq : in  std_logic                     := 'X'; -- irq
			receiver4_irq : in  std_logic                     := 'X'; -- irq
			receiver5_irq : in  std_logic                     := 'X'; -- irq
			receiver6_irq : in  std_logic                     := 'X'; -- irq
			receiver7_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component soc_system_v5_irq_mapper_001;

	component soc_system_v5_avalon_st_adapter is
		generic (
			inBitsPerSymbol : integer := 8;
			inUsePackets    : integer := 0;
			inDataWidth     : integer := 8;
			inChannelWidth  : integer := 3;
			inErrorWidth    : integer := 2;
			inUseEmptyPort  : integer := 0;
			inUseValid      : integer := 1;
			inUseReady      : integer := 1;
			inReadyLatency  : integer := 0;
			outDataWidth    : integer := 32;
			outChannelWidth : integer := 3;
			outErrorWidth   : integer := 2;
			outUseEmptyPort : integer := 0;
			outUseValid     : integer := 1;
			outUseReady     : integer := 1;
			outReadyLatency : integer := 0
		);
		port (
			in_clk_0_clk   : in  std_logic                     := 'X';             -- clk
			in_rst_0_reset : in  std_logic                     := 'X';             -- reset
			in_0_data      : in  std_logic_vector(15 downto 0) := (others => 'X'); -- data
			in_0_valid     : in  std_logic                     := 'X';             -- valid
			in_0_ready     : out std_logic;                                        -- ready
			out_0_data     : out std_logic_vector(31 downto 0);                    -- data
			out_0_valid    : out std_logic;                                        -- valid
			out_0_ready    : in  std_logic                     := 'X'              -- ready
		);
	end component soc_system_v5_avalon_st_adapter;

	component soc_system_v5_avalon_st_adapter_001 is
		generic (
			inBitsPerSymbol : integer := 8;
			inUsePackets    : integer := 0;
			inDataWidth     : integer := 8;
			inChannelWidth  : integer := 3;
			inErrorWidth    : integer := 2;
			inUseEmptyPort  : integer := 0;
			inUseValid      : integer := 1;
			inUseReady      : integer := 1;
			inReadyLatency  : integer := 0;
			outDataWidth    : integer := 32;
			outChannelWidth : integer := 3;
			outErrorWidth   : integer := 2;
			outUseEmptyPort : integer := 0;
			outUseValid     : integer := 1;
			outUseReady     : integer := 1;
			outReadyLatency : integer := 0
		);
		port (
			in_clk_0_clk   : in  std_logic                     := 'X';             -- clk
			in_rst_0_reset : in  std_logic                     := 'X';             -- reset
			in_0_data      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			in_0_valid     : in  std_logic                     := 'X';             -- valid
			in_0_ready     : out std_logic;                                        -- ready
			out_0_data     : out std_logic_vector(31 downto 0);                    -- data
			out_0_valid    : out std_logic;                                        -- valid
			out_0_ready    : in  std_logic                     := 'X'              -- ready
		);
	end component soc_system_v5_avalon_st_adapter_001;

	component soc_system_v5_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component soc_system_v5_rst_controller;

	component soc_system_v5_rst_controller_002 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component soc_system_v5_rst_controller_002;

	component soc_system_v5_adc_fifo_dc is
		generic (
			SYMBOLS_PER_BEAT   : integer := 1;
			BITS_PER_SYMBOL    : integer := 8;
			FIFO_DEPTH         : integer := 16;
			CHANNEL_WIDTH      : integer := 0;
			ERROR_WIDTH        : integer := 0;
			USE_PACKETS        : integer := 0;
			USE_IN_FILL_LEVEL  : integer := 0;
			USE_OUT_FILL_LEVEL : integer := 0;
			WR_SYNC_DEPTH      : integer := 3;
			RD_SYNC_DEPTH      : integer := 3
		);
		port (
			in_clk            : in  std_logic                     := 'X';             --        in_clk.clk
			in_reset_n        : in  std_logic                     := 'X';             --  in_clk_reset.reset_n
			out_clk           : in  std_logic                     := 'X';             --       out_clk.clk
			out_reset_n       : in  std_logic                     := 'X';             -- out_clk_reset.reset_n
			in_data           : in  std_logic_vector(15 downto 0) := (others => 'X'); --            in.data
			in_valid          : in  std_logic                     := 'X';             --              .valid
			in_ready          : out std_logic;                                        --              .ready
			out_data          : out std_logic_vector(15 downto 0);                    --           out.data
			out_valid         : out std_logic;                                        --              .valid
			out_ready         : in  std_logic                     := 'X';             --              .ready
			in_channel        : in  std_logic_vector(0 downto 0)  := (others => 'X');
			in_csr_address    : in  std_logic                     := 'X';
			in_csr_read       : in  std_logic                     := 'X';
			in_csr_readdata   : out std_logic_vector(31 downto 0);
			in_csr_write      : in  std_logic                     := 'X';
			in_csr_writedata  : in  std_logic_vector(31 downto 0) := (others => 'X');
			in_empty          : in  std_logic_vector(0 downto 0)  := (others => 'X');
			in_endofpacket    : in  std_logic                     := 'X';
			in_error          : in  std_logic_vector(0 downto 0)  := (others => 'X');
			in_startofpacket  : in  std_logic                     := 'X';
			out_channel       : out std_logic_vector(0 downto 0);
			out_csr_address   : in  std_logic                     := 'X';
			out_csr_read      : in  std_logic                     := 'X';
			out_csr_readdata  : out std_logic_vector(31 downto 0);
			out_csr_write     : in  std_logic                     := 'X';
			out_csr_writedata : in  std_logic_vector(31 downto 0) := (others => 'X');
			out_empty         : out std_logic_vector(0 downto 0);
			out_endofpacket   : out std_logic;
			out_error         : out std_logic_vector(0 downto 0);
			out_startofpacket : out std_logic;
			space_avail_data  : out std_logic_vector(14 downto 0)
		);
	end component soc_system_v5_adc_fifo_dc;

	component soc_system_v5_dconv_fifo_dc is
		generic (
			SYMBOLS_PER_BEAT   : integer := 1;
			BITS_PER_SYMBOL    : integer := 8;
			FIFO_DEPTH         : integer := 16;
			CHANNEL_WIDTH      : integer := 0;
			ERROR_WIDTH        : integer := 0;
			USE_PACKETS        : integer := 0;
			USE_IN_FILL_LEVEL  : integer := 0;
			USE_OUT_FILL_LEVEL : integer := 0;
			WR_SYNC_DEPTH      : integer := 3;
			RD_SYNC_DEPTH      : integer := 3
		);
		port (
			in_clk            : in  std_logic                     := 'X';             --        in_clk.clk
			in_reset_n        : in  std_logic                     := 'X';             --  in_clk_reset.reset_n
			out_clk           : in  std_logic                     := 'X';             --       out_clk.clk
			out_reset_n       : in  std_logic                     := 'X';             -- out_clk_reset.reset_n
			in_data           : in  std_logic_vector(31 downto 0) := (others => 'X'); --            in.data
			in_valid          : in  std_logic                     := 'X';             --              .valid
			in_ready          : out std_logic;                                        --              .ready
			out_data          : out std_logic_vector(31 downto 0);                    --           out.data
			out_valid         : out std_logic;                                        --              .valid
			out_ready         : in  std_logic                     := 'X';             --              .ready
			in_channel        : in  std_logic_vector(0 downto 0)  := (others => 'X');
			in_csr_address    : in  std_logic                     := 'X';
			in_csr_read       : in  std_logic                     := 'X';
			in_csr_readdata   : out std_logic_vector(31 downto 0);
			in_csr_write      : in  std_logic                     := 'X';
			in_csr_writedata  : in  std_logic_vector(31 downto 0) := (others => 'X');
			in_empty          : in  std_logic_vector(0 downto 0)  := (others => 'X');
			in_endofpacket    : in  std_logic                     := 'X';
			in_error          : in  std_logic_vector(0 downto 0)  := (others => 'X');
			in_startofpacket  : in  std_logic                     := 'X';
			out_channel       : out std_logic_vector(0 downto 0);
			out_csr_address   : in  std_logic                     := 'X';
			out_csr_read      : in  std_logic                     := 'X';
			out_csr_readdata  : out std_logic_vector(31 downto 0);
			out_csr_write     : in  std_logic                     := 'X';
			out_csr_writedata : in  std_logic_vector(31 downto 0) := (others => 'X');
			out_empty         : out std_logic_vector(0 downto 0);
			out_endofpacket   : out std_logic;
			out_error         : out std_logic_vector(0 downto 0);
			out_startofpacket : out std_logic;
			space_avail_data  : out std_logic_vector(15 downto 0)
		);
	end component soc_system_v5_dconv_fifo_dc;

	signal hps_0_h2f_reset_reset                                                 : std_logic;                      -- hps_0:h2f_rst_n -> [hps_0_h2f_reset_reset_n, hps_0_h2f_reset_reset_n:in]
	signal alt_vip_vfr_vga_avalon_streaming_source_valid                         : std_logic;                      -- alt_vip_vfr_vga:dout_valid -> alt_vip_itc_0:is_valid
	signal alt_vip_vfr_vga_avalon_streaming_source_data                          : std_logic_vector(31 downto 0);  -- alt_vip_vfr_vga:dout_data -> alt_vip_itc_0:is_data
	signal alt_vip_vfr_vga_avalon_streaming_source_ready                         : std_logic;                      -- alt_vip_itc_0:is_ready -> alt_vip_vfr_vga:dout_ready
	signal alt_vip_vfr_vga_avalon_streaming_source_startofpacket                 : std_logic;                      -- alt_vip_vfr_vga:dout_startofpacket -> alt_vip_itc_0:is_sop
	signal alt_vip_vfr_vga_avalon_streaming_source_endofpacket                   : std_logic;                      -- alt_vip_vfr_vga:dout_endofpacket -> alt_vip_itc_0:is_eop
	signal fifo_dummy64_in_out_valid                                             : std_logic;                      -- fifo_dummy64_in:avalonst_source_valid -> fifo_dummy64_out:avalonst_sink_valid
	signal fifo_dummy64_in_out_data                                              : std_logic_vector(31 downto 0);  -- fifo_dummy64_in:avalonst_source_data -> fifo_dummy64_out:avalonst_sink_data
	signal fifo_dummy64_in_out_ready                                             : std_logic;                      -- fifo_dummy64_out:avalonst_sink_ready -> fifo_dummy64_in:avalonst_source_ready
	signal gp_pll_outclk0_clk                                                    : std_logic;                      -- gp_pll:outclk_0 -> [alt_vip_itc_0:is_clk, alt_vip_vfr_vga:clock, mm_interconnect_1:gp_pll_outclk0_clk, rst_controller_002:clk]
	signal nmr_sys_pll_reconfig_from_pll_reconfig_from_pll                       : std_logic_vector(63 downto 0);  -- nmr_sys_pll:reconfig_from_pll -> nmr_sys_pll_reconfig:reconfig_from_pll
	signal analyzer_pll_reconfig_from_pll_reconfig_from_pll                      : std_logic_vector(63 downto 0);  -- analyzer_pll:reconfig_from_pll -> analyzer_pll_reconfig:reconfig_from_pll
	signal nmr_sys_pll_reconfig_reconfig_to_pll_reconfig_to_pll                  : std_logic_vector(63 downto 0);  -- nmr_sys_pll_reconfig:reconfig_to_pll -> nmr_sys_pll:reconfig_to_pll
	signal analyzer_pll_reconfig_reconfig_to_pll_reconfig_to_pll                 : std_logic_vector(63 downto 0);  -- analyzer_pll_reconfig:reconfig_to_pll -> analyzer_pll:reconfig_to_pll
	signal alt_vip_vfr_vga_avalon_master_readdata                                : std_logic_vector(127 downto 0); -- mm_interconnect_0:alt_vip_vfr_vga_avalon_master_readdata -> alt_vip_vfr_vga:master_readdata
	signal alt_vip_vfr_vga_avalon_master_waitrequest                             : std_logic;                      -- mm_interconnect_0:alt_vip_vfr_vga_avalon_master_waitrequest -> alt_vip_vfr_vga:master_waitrequest
	signal alt_vip_vfr_vga_avalon_master_address                                 : std_logic_vector(31 downto 0);  -- alt_vip_vfr_vga:master_address -> mm_interconnect_0:alt_vip_vfr_vga_avalon_master_address
	signal alt_vip_vfr_vga_avalon_master_read                                    : std_logic;                      -- alt_vip_vfr_vga:master_read -> mm_interconnect_0:alt_vip_vfr_vga_avalon_master_read
	signal alt_vip_vfr_vga_avalon_master_readdatavalid                           : std_logic;                      -- mm_interconnect_0:alt_vip_vfr_vga_avalon_master_readdatavalid -> alt_vip_vfr_vga:master_readdatavalid
	signal alt_vip_vfr_vga_avalon_master_burstcount                              : std_logic_vector(5 downto 0);   -- alt_vip_vfr_vga:master_burstcount -> mm_interconnect_0:alt_vip_vfr_vga_avalon_master_burstcount
	signal master_secure_master_readdata                                         : std_logic_vector(31 downto 0);  -- mm_interconnect_0:master_secure_master_readdata -> master_secure:master_readdata
	signal master_secure_master_waitrequest                                      : std_logic;                      -- mm_interconnect_0:master_secure_master_waitrequest -> master_secure:master_waitrequest
	signal master_secure_master_address                                          : std_logic_vector(31 downto 0);  -- master_secure:master_address -> mm_interconnect_0:master_secure_master_address
	signal master_secure_master_read                                             : std_logic;                      -- master_secure:master_read -> mm_interconnect_0:master_secure_master_read
	signal master_secure_master_byteenable                                       : std_logic_vector(3 downto 0);   -- master_secure:master_byteenable -> mm_interconnect_0:master_secure_master_byteenable
	signal master_secure_master_readdatavalid                                    : std_logic;                      -- mm_interconnect_0:master_secure_master_readdatavalid -> master_secure:master_readdatavalid
	signal master_secure_master_write                                            : std_logic;                      -- master_secure:master_write -> mm_interconnect_0:master_secure_master_write
	signal master_secure_master_writedata                                        : std_logic_vector(31 downto 0);  -- master_secure:master_writedata -> mm_interconnect_0:master_secure_master_writedata
	signal mm_interconnect_0_hps_0_f2h_axi_slave_awburst                         : std_logic_vector(1 downto 0);   -- mm_interconnect_0:hps_0_f2h_axi_slave_awburst -> hps_0:f2h_AWBURST
	signal mm_interconnect_0_hps_0_f2h_axi_slave_awuser                          : std_logic_vector(4 downto 0);   -- mm_interconnect_0:hps_0_f2h_axi_slave_awuser -> hps_0:f2h_AWUSER
	signal mm_interconnect_0_hps_0_f2h_axi_slave_arlen                           : std_logic_vector(3 downto 0);   -- mm_interconnect_0:hps_0_f2h_axi_slave_arlen -> hps_0:f2h_ARLEN
	signal mm_interconnect_0_hps_0_f2h_axi_slave_wstrb                           : std_logic_vector(15 downto 0);  -- mm_interconnect_0:hps_0_f2h_axi_slave_wstrb -> hps_0:f2h_WSTRB
	signal mm_interconnect_0_hps_0_f2h_axi_slave_wready                          : std_logic;                      -- hps_0:f2h_WREADY -> mm_interconnect_0:hps_0_f2h_axi_slave_wready
	signal mm_interconnect_0_hps_0_f2h_axi_slave_rid                             : std_logic_vector(7 downto 0);   -- hps_0:f2h_RID -> mm_interconnect_0:hps_0_f2h_axi_slave_rid
	signal mm_interconnect_0_hps_0_f2h_axi_slave_rready                          : std_logic;                      -- mm_interconnect_0:hps_0_f2h_axi_slave_rready -> hps_0:f2h_RREADY
	signal mm_interconnect_0_hps_0_f2h_axi_slave_awlen                           : std_logic_vector(3 downto 0);   -- mm_interconnect_0:hps_0_f2h_axi_slave_awlen -> hps_0:f2h_AWLEN
	signal mm_interconnect_0_hps_0_f2h_axi_slave_wid                             : std_logic_vector(7 downto 0);   -- mm_interconnect_0:hps_0_f2h_axi_slave_wid -> hps_0:f2h_WID
	signal mm_interconnect_0_hps_0_f2h_axi_slave_arcache                         : std_logic_vector(3 downto 0);   -- mm_interconnect_0:hps_0_f2h_axi_slave_arcache -> hps_0:f2h_ARCACHE
	signal mm_interconnect_0_hps_0_f2h_axi_slave_wvalid                          : std_logic;                      -- mm_interconnect_0:hps_0_f2h_axi_slave_wvalid -> hps_0:f2h_WVALID
	signal mm_interconnect_0_hps_0_f2h_axi_slave_araddr                          : std_logic_vector(31 downto 0);  -- mm_interconnect_0:hps_0_f2h_axi_slave_araddr -> hps_0:f2h_ARADDR
	signal mm_interconnect_0_hps_0_f2h_axi_slave_arprot                          : std_logic_vector(2 downto 0);   -- mm_interconnect_0:hps_0_f2h_axi_slave_arprot -> hps_0:f2h_ARPROT
	signal mm_interconnect_0_hps_0_f2h_axi_slave_awprot                          : std_logic_vector(2 downto 0);   -- mm_interconnect_0:hps_0_f2h_axi_slave_awprot -> hps_0:f2h_AWPROT
	signal mm_interconnect_0_hps_0_f2h_axi_slave_wdata                           : std_logic_vector(127 downto 0); -- mm_interconnect_0:hps_0_f2h_axi_slave_wdata -> hps_0:f2h_WDATA
	signal mm_interconnect_0_hps_0_f2h_axi_slave_arvalid                         : std_logic;                      -- mm_interconnect_0:hps_0_f2h_axi_slave_arvalid -> hps_0:f2h_ARVALID
	signal mm_interconnect_0_hps_0_f2h_axi_slave_awcache                         : std_logic_vector(3 downto 0);   -- mm_interconnect_0:hps_0_f2h_axi_slave_awcache -> hps_0:f2h_AWCACHE
	signal mm_interconnect_0_hps_0_f2h_axi_slave_arid                            : std_logic_vector(7 downto 0);   -- mm_interconnect_0:hps_0_f2h_axi_slave_arid -> hps_0:f2h_ARID
	signal mm_interconnect_0_hps_0_f2h_axi_slave_arlock                          : std_logic_vector(1 downto 0);   -- mm_interconnect_0:hps_0_f2h_axi_slave_arlock -> hps_0:f2h_ARLOCK
	signal mm_interconnect_0_hps_0_f2h_axi_slave_awlock                          : std_logic_vector(1 downto 0);   -- mm_interconnect_0:hps_0_f2h_axi_slave_awlock -> hps_0:f2h_AWLOCK
	signal mm_interconnect_0_hps_0_f2h_axi_slave_awaddr                          : std_logic_vector(31 downto 0);  -- mm_interconnect_0:hps_0_f2h_axi_slave_awaddr -> hps_0:f2h_AWADDR
	signal mm_interconnect_0_hps_0_f2h_axi_slave_bresp                           : std_logic_vector(1 downto 0);   -- hps_0:f2h_BRESP -> mm_interconnect_0:hps_0_f2h_axi_slave_bresp
	signal mm_interconnect_0_hps_0_f2h_axi_slave_arready                         : std_logic;                      -- hps_0:f2h_ARREADY -> mm_interconnect_0:hps_0_f2h_axi_slave_arready
	signal mm_interconnect_0_hps_0_f2h_axi_slave_rdata                           : std_logic_vector(127 downto 0); -- hps_0:f2h_RDATA -> mm_interconnect_0:hps_0_f2h_axi_slave_rdata
	signal mm_interconnect_0_hps_0_f2h_axi_slave_awready                         : std_logic;                      -- hps_0:f2h_AWREADY -> mm_interconnect_0:hps_0_f2h_axi_slave_awready
	signal mm_interconnect_0_hps_0_f2h_axi_slave_arburst                         : std_logic_vector(1 downto 0);   -- mm_interconnect_0:hps_0_f2h_axi_slave_arburst -> hps_0:f2h_ARBURST
	signal mm_interconnect_0_hps_0_f2h_axi_slave_arsize                          : std_logic_vector(2 downto 0);   -- mm_interconnect_0:hps_0_f2h_axi_slave_arsize -> hps_0:f2h_ARSIZE
	signal mm_interconnect_0_hps_0_f2h_axi_slave_bready                          : std_logic;                      -- mm_interconnect_0:hps_0_f2h_axi_slave_bready -> hps_0:f2h_BREADY
	signal mm_interconnect_0_hps_0_f2h_axi_slave_rlast                           : std_logic;                      -- hps_0:f2h_RLAST -> mm_interconnect_0:hps_0_f2h_axi_slave_rlast
	signal mm_interconnect_0_hps_0_f2h_axi_slave_wlast                           : std_logic;                      -- mm_interconnect_0:hps_0_f2h_axi_slave_wlast -> hps_0:f2h_WLAST
	signal mm_interconnect_0_hps_0_f2h_axi_slave_rresp                           : std_logic_vector(1 downto 0);   -- hps_0:f2h_RRESP -> mm_interconnect_0:hps_0_f2h_axi_slave_rresp
	signal mm_interconnect_0_hps_0_f2h_axi_slave_awid                            : std_logic_vector(7 downto 0);   -- mm_interconnect_0:hps_0_f2h_axi_slave_awid -> hps_0:f2h_AWID
	signal mm_interconnect_0_hps_0_f2h_axi_slave_bid                             : std_logic_vector(7 downto 0);   -- hps_0:f2h_BID -> mm_interconnect_0:hps_0_f2h_axi_slave_bid
	signal mm_interconnect_0_hps_0_f2h_axi_slave_bvalid                          : std_logic;                      -- hps_0:f2h_BVALID -> mm_interconnect_0:hps_0_f2h_axi_slave_bvalid
	signal mm_interconnect_0_hps_0_f2h_axi_slave_awsize                          : std_logic_vector(2 downto 0);   -- mm_interconnect_0:hps_0_f2h_axi_slave_awsize -> hps_0:f2h_AWSIZE
	signal mm_interconnect_0_hps_0_f2h_axi_slave_awvalid                         : std_logic;                      -- mm_interconnect_0:hps_0_f2h_axi_slave_awvalid -> hps_0:f2h_AWVALID
	signal mm_interconnect_0_hps_0_f2h_axi_slave_aruser                          : std_logic_vector(4 downto 0);   -- mm_interconnect_0:hps_0_f2h_axi_slave_aruser -> hps_0:f2h_ARUSER
	signal mm_interconnect_0_hps_0_f2h_axi_slave_rvalid                          : std_logic;                      -- hps_0:f2h_RVALID -> mm_interconnect_0:hps_0_f2h_axi_slave_rvalid
	signal hps_0_h2f_axi_master_awburst                                          : std_logic_vector(1 downto 0);   -- hps_0:h2f_AWBURST -> mm_interconnect_1:hps_0_h2f_axi_master_awburst
	signal hps_0_h2f_axi_master_arlen                                            : std_logic_vector(3 downto 0);   -- hps_0:h2f_ARLEN -> mm_interconnect_1:hps_0_h2f_axi_master_arlen
	signal hps_0_h2f_axi_master_wstrb                                            : std_logic_vector(15 downto 0);  -- hps_0:h2f_WSTRB -> mm_interconnect_1:hps_0_h2f_axi_master_wstrb
	signal hps_0_h2f_axi_master_wready                                           : std_logic;                      -- mm_interconnect_1:hps_0_h2f_axi_master_wready -> hps_0:h2f_WREADY
	signal hps_0_h2f_axi_master_rid                                              : std_logic_vector(11 downto 0);  -- mm_interconnect_1:hps_0_h2f_axi_master_rid -> hps_0:h2f_RID
	signal hps_0_h2f_axi_master_rready                                           : std_logic;                      -- hps_0:h2f_RREADY -> mm_interconnect_1:hps_0_h2f_axi_master_rready
	signal hps_0_h2f_axi_master_awlen                                            : std_logic_vector(3 downto 0);   -- hps_0:h2f_AWLEN -> mm_interconnect_1:hps_0_h2f_axi_master_awlen
	signal hps_0_h2f_axi_master_wid                                              : std_logic_vector(11 downto 0);  -- hps_0:h2f_WID -> mm_interconnect_1:hps_0_h2f_axi_master_wid
	signal hps_0_h2f_axi_master_arcache                                          : std_logic_vector(3 downto 0);   -- hps_0:h2f_ARCACHE -> mm_interconnect_1:hps_0_h2f_axi_master_arcache
	signal hps_0_h2f_axi_master_wvalid                                           : std_logic;                      -- hps_0:h2f_WVALID -> mm_interconnect_1:hps_0_h2f_axi_master_wvalid
	signal hps_0_h2f_axi_master_araddr                                           : std_logic_vector(29 downto 0);  -- hps_0:h2f_ARADDR -> mm_interconnect_1:hps_0_h2f_axi_master_araddr
	signal hps_0_h2f_axi_master_arprot                                           : std_logic_vector(2 downto 0);   -- hps_0:h2f_ARPROT -> mm_interconnect_1:hps_0_h2f_axi_master_arprot
	signal hps_0_h2f_axi_master_awprot                                           : std_logic_vector(2 downto 0);   -- hps_0:h2f_AWPROT -> mm_interconnect_1:hps_0_h2f_axi_master_awprot
	signal hps_0_h2f_axi_master_wdata                                            : std_logic_vector(127 downto 0); -- hps_0:h2f_WDATA -> mm_interconnect_1:hps_0_h2f_axi_master_wdata
	signal hps_0_h2f_axi_master_arvalid                                          : std_logic;                      -- hps_0:h2f_ARVALID -> mm_interconnect_1:hps_0_h2f_axi_master_arvalid
	signal hps_0_h2f_axi_master_awcache                                          : std_logic_vector(3 downto 0);   -- hps_0:h2f_AWCACHE -> mm_interconnect_1:hps_0_h2f_axi_master_awcache
	signal hps_0_h2f_axi_master_arid                                             : std_logic_vector(11 downto 0);  -- hps_0:h2f_ARID -> mm_interconnect_1:hps_0_h2f_axi_master_arid
	signal hps_0_h2f_axi_master_arlock                                           : std_logic_vector(1 downto 0);   -- hps_0:h2f_ARLOCK -> mm_interconnect_1:hps_0_h2f_axi_master_arlock
	signal hps_0_h2f_axi_master_awlock                                           : std_logic_vector(1 downto 0);   -- hps_0:h2f_AWLOCK -> mm_interconnect_1:hps_0_h2f_axi_master_awlock
	signal hps_0_h2f_axi_master_awaddr                                           : std_logic_vector(29 downto 0);  -- hps_0:h2f_AWADDR -> mm_interconnect_1:hps_0_h2f_axi_master_awaddr
	signal hps_0_h2f_axi_master_bresp                                            : std_logic_vector(1 downto 0);   -- mm_interconnect_1:hps_0_h2f_axi_master_bresp -> hps_0:h2f_BRESP
	signal hps_0_h2f_axi_master_arready                                          : std_logic;                      -- mm_interconnect_1:hps_0_h2f_axi_master_arready -> hps_0:h2f_ARREADY
	signal hps_0_h2f_axi_master_rdata                                            : std_logic_vector(127 downto 0); -- mm_interconnect_1:hps_0_h2f_axi_master_rdata -> hps_0:h2f_RDATA
	signal hps_0_h2f_axi_master_awready                                          : std_logic;                      -- mm_interconnect_1:hps_0_h2f_axi_master_awready -> hps_0:h2f_AWREADY
	signal hps_0_h2f_axi_master_arburst                                          : std_logic_vector(1 downto 0);   -- hps_0:h2f_ARBURST -> mm_interconnect_1:hps_0_h2f_axi_master_arburst
	signal hps_0_h2f_axi_master_arsize                                           : std_logic_vector(2 downto 0);   -- hps_0:h2f_ARSIZE -> mm_interconnect_1:hps_0_h2f_axi_master_arsize
	signal hps_0_h2f_axi_master_bready                                           : std_logic;                      -- hps_0:h2f_BREADY -> mm_interconnect_1:hps_0_h2f_axi_master_bready
	signal hps_0_h2f_axi_master_rlast                                            : std_logic;                      -- mm_interconnect_1:hps_0_h2f_axi_master_rlast -> hps_0:h2f_RLAST
	signal hps_0_h2f_axi_master_wlast                                            : std_logic;                      -- hps_0:h2f_WLAST -> mm_interconnect_1:hps_0_h2f_axi_master_wlast
	signal hps_0_h2f_axi_master_rresp                                            : std_logic_vector(1 downto 0);   -- mm_interconnect_1:hps_0_h2f_axi_master_rresp -> hps_0:h2f_RRESP
	signal hps_0_h2f_axi_master_awid                                             : std_logic_vector(11 downto 0);  -- hps_0:h2f_AWID -> mm_interconnect_1:hps_0_h2f_axi_master_awid
	signal hps_0_h2f_axi_master_bid                                              : std_logic_vector(11 downto 0);  -- mm_interconnect_1:hps_0_h2f_axi_master_bid -> hps_0:h2f_BID
	signal hps_0_h2f_axi_master_bvalid                                           : std_logic;                      -- mm_interconnect_1:hps_0_h2f_axi_master_bvalid -> hps_0:h2f_BVALID
	signal hps_0_h2f_axi_master_awsize                                           : std_logic_vector(2 downto 0);   -- hps_0:h2f_AWSIZE -> mm_interconnect_1:hps_0_h2f_axi_master_awsize
	signal hps_0_h2f_axi_master_awvalid                                          : std_logic;                      -- hps_0:h2f_AWVALID -> mm_interconnect_1:hps_0_h2f_axi_master_awvalid
	signal hps_0_h2f_axi_master_rvalid                                           : std_logic;                      -- mm_interconnect_1:hps_0_h2f_axi_master_rvalid -> hps_0:h2f_RVALID
	signal dma_fifo_write_master_chipselect                                      : std_logic;                      -- dma_fifo:write_chipselect -> mm_interconnect_1:dma_fifo_write_master_chipselect
	signal dma_fifo_write_master_waitrequest                                     : std_logic;                      -- mm_interconnect_1:dma_fifo_write_master_waitrequest -> dma_fifo:write_waitrequest
	signal dma_fifo_write_master_address                                         : std_logic_vector(25 downto 0);  -- dma_fifo:write_address -> mm_interconnect_1:dma_fifo_write_master_address
	signal dma_fifo_write_master_byteenable                                      : std_logic_vector(3 downto 0);   -- dma_fifo:write_byteenable -> mm_interconnect_1:dma_fifo_write_master_byteenable
	signal dma_fifo_write_master_write                                           : std_logic;                      -- dma_fifo:write_write_n -> dma_fifo_write_master_write:in
	signal dma_fifo_write_master_writedata                                       : std_logic_vector(31 downto 0);  -- dma_fifo:write_writedata -> mm_interconnect_1:dma_fifo_write_master_writedata
	signal dma_dconvi_write_master_chipselect                                    : std_logic;                      -- dma_dconvi:write_chipselect -> mm_interconnect_1:dma_dconvi_write_master_chipselect
	signal dma_dconvi_write_master_waitrequest                                   : std_logic;                      -- mm_interconnect_1:dma_dconvi_write_master_waitrequest -> dma_dconvi:write_waitrequest
	signal dma_dconvi_write_master_address                                       : std_logic_vector(25 downto 0);  -- dma_dconvi:write_address -> mm_interconnect_1:dma_dconvi_write_master_address
	signal dma_dconvi_write_master_byteenable                                    : std_logic_vector(3 downto 0);   -- dma_dconvi:write_byteenable -> mm_interconnect_1:dma_dconvi_write_master_byteenable
	signal dma_dconvi_write_master_write                                         : std_logic;                      -- dma_dconvi:write_write_n -> dma_dconvi_write_master_write:in
	signal dma_dconvi_write_master_writedata                                     : std_logic_vector(31 downto 0);  -- dma_dconvi:write_writedata -> mm_interconnect_1:dma_dconvi_write_master_writedata
	signal dma_dconvq_write_master_chipselect                                    : std_logic;                      -- dma_dconvq:write_chipselect -> mm_interconnect_1:dma_dconvq_write_master_chipselect
	signal dma_dconvq_write_master_waitrequest                                   : std_logic;                      -- mm_interconnect_1:dma_dconvq_write_master_waitrequest -> dma_dconvq:write_waitrequest
	signal dma_dconvq_write_master_address                                       : std_logic_vector(25 downto 0);  -- dma_dconvq:write_address -> mm_interconnect_1:dma_dconvq_write_master_address
	signal dma_dconvq_write_master_byteenable                                    : std_logic_vector(3 downto 0);   -- dma_dconvq:write_byteenable -> mm_interconnect_1:dma_dconvq_write_master_byteenable
	signal dma_dconvq_write_master_write                                         : std_logic;                      -- dma_dconvq:write_write_n -> dma_dconvq_write_master_write:in
	signal dma_dconvq_write_master_writedata                                     : std_logic_vector(31 downto 0);  -- dma_dconvq:write_writedata -> mm_interconnect_1:dma_dconvq_write_master_writedata
	signal dma_dummy_write_master_chipselect                                     : std_logic;                      -- dma_dummy:write_chipselect -> mm_interconnect_1:dma_dummy_write_master_chipselect
	signal dma_dummy_write_master_waitrequest                                    : std_logic;                      -- mm_interconnect_1:dma_dummy_write_master_waitrequest -> dma_dummy:write_waitrequest
	signal dma_dummy_write_master_address                                        : std_logic_vector(25 downto 0);  -- dma_dummy:write_address -> mm_interconnect_1:dma_dummy_write_master_address
	signal dma_dummy_write_master_byteenable                                     : std_logic_vector(3 downto 0);   -- dma_dummy:write_byteenable -> mm_interconnect_1:dma_dummy_write_master_byteenable
	signal dma_dummy_write_master_write                                          : std_logic;                      -- dma_dummy:write_write_n -> dma_dummy_write_master_write:in
	signal dma_dummy_write_master_writedata                                      : std_logic_vector(31 downto 0);  -- dma_dummy:write_writedata -> mm_interconnect_1:dma_dummy_write_master_writedata
	signal dma_fifo_read_master_chipselect                                       : std_logic;                      -- dma_fifo:read_chipselect -> mm_interconnect_1:dma_fifo_read_master_chipselect
	signal dma_fifo_read_master_readdata                                         : std_logic_vector(31 downto 0);  -- mm_interconnect_1:dma_fifo_read_master_readdata -> dma_fifo:read_readdata
	signal dma_fifo_read_master_waitrequest                                      : std_logic;                      -- mm_interconnect_1:dma_fifo_read_master_waitrequest -> dma_fifo:read_waitrequest
	signal dma_fifo_read_master_address                                          : std_logic_vector(26 downto 0);  -- dma_fifo:read_address -> mm_interconnect_1:dma_fifo_read_master_address
	signal dma_fifo_read_master_read                                             : std_logic;                      -- dma_fifo:read_read_n -> dma_fifo_read_master_read:in
	signal dma_fifo_read_master_readdatavalid                                    : std_logic;                      -- mm_interconnect_1:dma_fifo_read_master_readdatavalid -> dma_fifo:read_readdatavalid
	signal hps_0_h2f_lw_axi_master_awburst                                       : std_logic_vector(1 downto 0);   -- hps_0:h2f_lw_AWBURST -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awburst
	signal hps_0_h2f_lw_axi_master_arlen                                         : std_logic_vector(3 downto 0);   -- hps_0:h2f_lw_ARLEN -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arlen
	signal hps_0_h2f_lw_axi_master_wstrb                                         : std_logic_vector(3 downto 0);   -- hps_0:h2f_lw_WSTRB -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wstrb
	signal hps_0_h2f_lw_axi_master_wready                                        : std_logic;                      -- mm_interconnect_1:hps_0_h2f_lw_axi_master_wready -> hps_0:h2f_lw_WREADY
	signal hps_0_h2f_lw_axi_master_rid                                           : std_logic_vector(11 downto 0);  -- mm_interconnect_1:hps_0_h2f_lw_axi_master_rid -> hps_0:h2f_lw_RID
	signal hps_0_h2f_lw_axi_master_rready                                        : std_logic;                      -- hps_0:h2f_lw_RREADY -> mm_interconnect_1:hps_0_h2f_lw_axi_master_rready
	signal hps_0_h2f_lw_axi_master_awlen                                         : std_logic_vector(3 downto 0);   -- hps_0:h2f_lw_AWLEN -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awlen
	signal hps_0_h2f_lw_axi_master_wid                                           : std_logic_vector(11 downto 0);  -- hps_0:h2f_lw_WID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wid
	signal hps_0_h2f_lw_axi_master_arcache                                       : std_logic_vector(3 downto 0);   -- hps_0:h2f_lw_ARCACHE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arcache
	signal hps_0_h2f_lw_axi_master_wvalid                                        : std_logic;                      -- hps_0:h2f_lw_WVALID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wvalid
	signal hps_0_h2f_lw_axi_master_araddr                                        : std_logic_vector(20 downto 0);  -- hps_0:h2f_lw_ARADDR -> mm_interconnect_1:hps_0_h2f_lw_axi_master_araddr
	signal hps_0_h2f_lw_axi_master_arprot                                        : std_logic_vector(2 downto 0);   -- hps_0:h2f_lw_ARPROT -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arprot
	signal hps_0_h2f_lw_axi_master_awprot                                        : std_logic_vector(2 downto 0);   -- hps_0:h2f_lw_AWPROT -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awprot
	signal hps_0_h2f_lw_axi_master_wdata                                         : std_logic_vector(31 downto 0);  -- hps_0:h2f_lw_WDATA -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wdata
	signal hps_0_h2f_lw_axi_master_arvalid                                       : std_logic;                      -- hps_0:h2f_lw_ARVALID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arvalid
	signal hps_0_h2f_lw_axi_master_awcache                                       : std_logic_vector(3 downto 0);   -- hps_0:h2f_lw_AWCACHE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awcache
	signal hps_0_h2f_lw_axi_master_arid                                          : std_logic_vector(11 downto 0);  -- hps_0:h2f_lw_ARID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arid
	signal hps_0_h2f_lw_axi_master_arlock                                        : std_logic_vector(1 downto 0);   -- hps_0:h2f_lw_ARLOCK -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arlock
	signal hps_0_h2f_lw_axi_master_awlock                                        : std_logic_vector(1 downto 0);   -- hps_0:h2f_lw_AWLOCK -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awlock
	signal hps_0_h2f_lw_axi_master_awaddr                                        : std_logic_vector(20 downto 0);  -- hps_0:h2f_lw_AWADDR -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awaddr
	signal hps_0_h2f_lw_axi_master_bresp                                         : std_logic_vector(1 downto 0);   -- mm_interconnect_1:hps_0_h2f_lw_axi_master_bresp -> hps_0:h2f_lw_BRESP
	signal hps_0_h2f_lw_axi_master_arready                                       : std_logic;                      -- mm_interconnect_1:hps_0_h2f_lw_axi_master_arready -> hps_0:h2f_lw_ARREADY
	signal hps_0_h2f_lw_axi_master_rdata                                         : std_logic_vector(31 downto 0);  -- mm_interconnect_1:hps_0_h2f_lw_axi_master_rdata -> hps_0:h2f_lw_RDATA
	signal hps_0_h2f_lw_axi_master_awready                                       : std_logic;                      -- mm_interconnect_1:hps_0_h2f_lw_axi_master_awready -> hps_0:h2f_lw_AWREADY
	signal hps_0_h2f_lw_axi_master_arburst                                       : std_logic_vector(1 downto 0);   -- hps_0:h2f_lw_ARBURST -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arburst
	signal hps_0_h2f_lw_axi_master_arsize                                        : std_logic_vector(2 downto 0);   -- hps_0:h2f_lw_ARSIZE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_arsize
	signal hps_0_h2f_lw_axi_master_bready                                        : std_logic;                      -- hps_0:h2f_lw_BREADY -> mm_interconnect_1:hps_0_h2f_lw_axi_master_bready
	signal hps_0_h2f_lw_axi_master_rlast                                         : std_logic;                      -- mm_interconnect_1:hps_0_h2f_lw_axi_master_rlast -> hps_0:h2f_lw_RLAST
	signal hps_0_h2f_lw_axi_master_wlast                                         : std_logic;                      -- hps_0:h2f_lw_WLAST -> mm_interconnect_1:hps_0_h2f_lw_axi_master_wlast
	signal hps_0_h2f_lw_axi_master_rresp                                         : std_logic_vector(1 downto 0);   -- mm_interconnect_1:hps_0_h2f_lw_axi_master_rresp -> hps_0:h2f_lw_RRESP
	signal hps_0_h2f_lw_axi_master_awid                                          : std_logic_vector(11 downto 0);  -- hps_0:h2f_lw_AWID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awid
	signal hps_0_h2f_lw_axi_master_bid                                           : std_logic_vector(11 downto 0);  -- mm_interconnect_1:hps_0_h2f_lw_axi_master_bid -> hps_0:h2f_lw_BID
	signal hps_0_h2f_lw_axi_master_bvalid                                        : std_logic;                      -- mm_interconnect_1:hps_0_h2f_lw_axi_master_bvalid -> hps_0:h2f_lw_BVALID
	signal hps_0_h2f_lw_axi_master_awsize                                        : std_logic_vector(2 downto 0);   -- hps_0:h2f_lw_AWSIZE -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awsize
	signal hps_0_h2f_lw_axi_master_awvalid                                       : std_logic;                      -- hps_0:h2f_lw_AWVALID -> mm_interconnect_1:hps_0_h2f_lw_axi_master_awvalid
	signal hps_0_h2f_lw_axi_master_rvalid                                        : std_logic;                      -- mm_interconnect_1:hps_0_h2f_lw_axi_master_rvalid -> hps_0:h2f_lw_RVALID
	signal master_non_sec_master_readdata                                        : std_logic_vector(31 downto 0);  -- mm_interconnect_1:master_non_sec_master_readdata -> master_non_sec:master_readdata
	signal master_non_sec_master_waitrequest                                     : std_logic;                      -- mm_interconnect_1:master_non_sec_master_waitrequest -> master_non_sec:master_waitrequest
	signal master_non_sec_master_address                                         : std_logic_vector(31 downto 0);  -- master_non_sec:master_address -> mm_interconnect_1:master_non_sec_master_address
	signal master_non_sec_master_read                                            : std_logic;                      -- master_non_sec:master_read -> mm_interconnect_1:master_non_sec_master_read
	signal master_non_sec_master_byteenable                                      : std_logic_vector(3 downto 0);   -- master_non_sec:master_byteenable -> mm_interconnect_1:master_non_sec_master_byteenable
	signal master_non_sec_master_readdatavalid                                   : std_logic;                      -- mm_interconnect_1:master_non_sec_master_readdatavalid -> master_non_sec:master_readdatavalid
	signal master_non_sec_master_write                                           : std_logic;                      -- master_non_sec:master_write -> mm_interconnect_1:master_non_sec_master_write
	signal master_non_sec_master_writedata                                       : std_logic_vector(31 downto 0);  -- master_non_sec:master_writedata -> mm_interconnect_1:master_non_sec_master_writedata
	signal dma_dconvq_read_master_chipselect                                     : std_logic;                      -- dma_dconvq:read_chipselect -> mm_interconnect_1:dma_dconvq_read_master_chipselect
	signal dma_dconvq_read_master_readdata                                       : std_logic_vector(31 downto 0);  -- mm_interconnect_1:dma_dconvq_read_master_readdata -> dma_dconvq:read_readdata
	signal dma_dconvq_read_master_waitrequest                                    : std_logic;                      -- mm_interconnect_1:dma_dconvq_read_master_waitrequest -> dma_dconvq:read_waitrequest
	signal dma_dconvq_read_master_address                                        : std_logic_vector(10 downto 0);  -- dma_dconvq:read_address -> mm_interconnect_1:dma_dconvq_read_master_address
	signal dma_dconvq_read_master_read                                           : std_logic;                      -- dma_dconvq:read_read_n -> dma_dconvq_read_master_read:in
	signal dma_dconvq_read_master_readdatavalid                                  : std_logic;                      -- mm_interconnect_1:dma_dconvq_read_master_readdatavalid -> dma_dconvq:read_readdatavalid
	signal dma_dconvi_read_master_chipselect                                     : std_logic;                      -- dma_dconvi:read_chipselect -> mm_interconnect_1:dma_dconvi_read_master_chipselect
	signal dma_dconvi_read_master_readdata                                       : std_logic_vector(31 downto 0);  -- mm_interconnect_1:dma_dconvi_read_master_readdata -> dma_dconvi:read_readdata
	signal dma_dconvi_read_master_waitrequest                                    : std_logic;                      -- mm_interconnect_1:dma_dconvi_read_master_waitrequest -> dma_dconvi:read_waitrequest
	signal dma_dconvi_read_master_address                                        : std_logic_vector(10 downto 0);  -- dma_dconvi:read_address -> mm_interconnect_1:dma_dconvi_read_master_address
	signal dma_dconvi_read_master_read                                           : std_logic;                      -- dma_dconvi:read_read_n -> dma_dconvi_read_master_read:in
	signal dma_dconvi_read_master_readdatavalid                                  : std_logic;                      -- mm_interconnect_1:dma_dconvi_read_master_readdatavalid -> dma_dconvi:read_readdatavalid
	signal dma_dummy_read_master_chipselect                                      : std_logic;                      -- dma_dummy:read_chipselect -> mm_interconnect_1:dma_dummy_read_master_chipselect
	signal dma_dummy_read_master_readdata                                        : std_logic_vector(31 downto 0);  -- mm_interconnect_1:dma_dummy_read_master_readdata -> dma_dummy:read_readdata
	signal dma_dummy_read_master_waitrequest                                     : std_logic;                      -- mm_interconnect_1:dma_dummy_read_master_waitrequest -> dma_dummy:read_waitrequest
	signal dma_dummy_read_master_address                                         : std_logic_vector(26 downto 0);  -- dma_dummy:read_address -> mm_interconnect_1:dma_dummy_read_master_address
	signal dma_dummy_read_master_read                                            : std_logic;                      -- dma_dummy:read_read_n -> dma_dummy_read_master_read:in
	signal dma_dummy_read_master_readdatavalid                                   : std_logic;                      -- mm_interconnect_1:dma_dummy_read_master_readdatavalid -> dma_dummy:read_readdatavalid
	signal mm_interconnect_1_fifo_dummy64_in_in_waitrequest                      : std_logic;                      -- fifo_dummy64_in:avalonmm_write_slave_waitrequest -> mm_interconnect_1:fifo_dummy64_in_in_waitrequest
	signal mm_interconnect_1_fifo_dummy64_in_in_address                          : std_logic_vector(0 downto 0);   -- mm_interconnect_1:fifo_dummy64_in_in_address -> fifo_dummy64_in:avalonmm_write_slave_address
	signal mm_interconnect_1_fifo_dummy64_in_in_write                            : std_logic;                      -- mm_interconnect_1:fifo_dummy64_in_in_write -> fifo_dummy64_in:avalonmm_write_slave_write
	signal mm_interconnect_1_fifo_dummy64_in_in_writedata                        : std_logic_vector(31 downto 0);  -- mm_interconnect_1:fifo_dummy64_in_in_writedata -> fifo_dummy64_in:avalonmm_write_slave_writedata
	signal mm_interconnect_1_fifo_dummy_in_waitrequest                           : std_logic;                      -- fifo_dummy:avalonmm_write_slave_waitrequest -> mm_interconnect_1:fifo_dummy_in_waitrequest
	signal mm_interconnect_1_fifo_dummy_in_write                                 : std_logic;                      -- mm_interconnect_1:fifo_dummy_in_write -> fifo_dummy:avalonmm_write_slave_write
	signal mm_interconnect_1_fifo_dummy_in_writedata                             : std_logic_vector(31 downto 0);  -- mm_interconnect_1:fifo_dummy_in_writedata -> fifo_dummy:avalonmm_write_slave_writedata
	signal mm_interconnect_1_fifo_dummy64_in_in_csr_readdata                     : std_logic_vector(31 downto 0);  -- fifo_dummy64_in:wrclk_control_slave_readdata -> mm_interconnect_1:fifo_dummy64_in_in_csr_readdata
	signal mm_interconnect_1_fifo_dummy64_in_in_csr_address                      : std_logic_vector(2 downto 0);   -- mm_interconnect_1:fifo_dummy64_in_in_csr_address -> fifo_dummy64_in:wrclk_control_slave_address
	signal mm_interconnect_1_fifo_dummy64_in_in_csr_read                         : std_logic;                      -- mm_interconnect_1:fifo_dummy64_in_in_csr_read -> fifo_dummy64_in:wrclk_control_slave_read
	signal mm_interconnect_1_fifo_dummy64_in_in_csr_write                        : std_logic;                      -- mm_interconnect_1:fifo_dummy64_in_in_csr_write -> fifo_dummy64_in:wrclk_control_slave_write
	signal mm_interconnect_1_fifo_dummy64_in_in_csr_writedata                    : std_logic_vector(31 downto 0);  -- mm_interconnect_1:fifo_dummy64_in_in_csr_writedata -> fifo_dummy64_in:wrclk_control_slave_writedata
	signal mm_interconnect_1_fifo_dummy64_out_in_csr_readdata                    : std_logic_vector(31 downto 0);  -- fifo_dummy64_out:wrclk_control_slave_readdata -> mm_interconnect_1:fifo_dummy64_out_in_csr_readdata
	signal mm_interconnect_1_fifo_dummy64_out_in_csr_address                     : std_logic_vector(2 downto 0);   -- mm_interconnect_1:fifo_dummy64_out_in_csr_address -> fifo_dummy64_out:wrclk_control_slave_address
	signal mm_interconnect_1_fifo_dummy64_out_in_csr_read                        : std_logic;                      -- mm_interconnect_1:fifo_dummy64_out_in_csr_read -> fifo_dummy64_out:wrclk_control_slave_read
	signal mm_interconnect_1_fifo_dummy64_out_in_csr_write                       : std_logic;                      -- mm_interconnect_1:fifo_dummy64_out_in_csr_write -> fifo_dummy64_out:wrclk_control_slave_write
	signal mm_interconnect_1_fifo_dummy64_out_in_csr_writedata                   : std_logic_vector(31 downto 0);  -- mm_interconnect_1:fifo_dummy64_out_in_csr_writedata -> fifo_dummy64_out:wrclk_control_slave_writedata
	signal mm_interconnect_1_fifo_dummy_in_csr_readdata                          : std_logic_vector(31 downto 0);  -- fifo_dummy:wrclk_control_slave_readdata -> mm_interconnect_1:fifo_dummy_in_csr_readdata
	signal mm_interconnect_1_fifo_dummy_in_csr_address                           : std_logic_vector(2 downto 0);   -- mm_interconnect_1:fifo_dummy_in_csr_address -> fifo_dummy:wrclk_control_slave_address
	signal mm_interconnect_1_fifo_dummy_in_csr_read                              : std_logic;                      -- mm_interconnect_1:fifo_dummy_in_csr_read -> fifo_dummy:wrclk_control_slave_read
	signal mm_interconnect_1_fifo_dummy_in_csr_write                             : std_logic;                      -- mm_interconnect_1:fifo_dummy_in_csr_write -> fifo_dummy:wrclk_control_slave_write
	signal mm_interconnect_1_fifo_dummy_in_csr_writedata                         : std_logic_vector(31 downto 0);  -- mm_interconnect_1:fifo_dummy_in_csr_writedata -> fifo_dummy:wrclk_control_slave_writedata
	signal mm_interconnect_1_fifo_dummy64_out_out_readdata                       : std_logic_vector(31 downto 0);  -- fifo_dummy64_out:avalonmm_read_slave_readdata -> mm_interconnect_1:fifo_dummy64_out_out_readdata
	signal mm_interconnect_1_fifo_dummy64_out_out_waitrequest                    : std_logic;                      -- fifo_dummy64_out:avalonmm_read_slave_waitrequest -> mm_interconnect_1:fifo_dummy64_out_out_waitrequest
	signal mm_interconnect_1_fifo_dummy64_out_out_address                        : std_logic_vector(0 downto 0);   -- mm_interconnect_1:fifo_dummy64_out_out_address -> fifo_dummy64_out:avalonmm_read_slave_address
	signal mm_interconnect_1_fifo_dummy64_out_out_read                           : std_logic;                      -- mm_interconnect_1:fifo_dummy64_out_out_read -> fifo_dummy64_out:avalonmm_read_slave_read
	signal mm_interconnect_1_fifo_dummy_out_readdata                             : std_logic_vector(31 downto 0);  -- fifo_dummy:avalonmm_read_slave_readdata -> mm_interconnect_1:fifo_dummy_out_readdata
	signal mm_interconnect_1_fifo_dummy_out_waitrequest                          : std_logic;                      -- fifo_dummy:avalonmm_read_slave_waitrequest -> mm_interconnect_1:fifo_dummy_out_waitrequest
	signal mm_interconnect_1_fifo_dummy_out_read                                 : std_logic;                      -- mm_interconnect_1:fifo_dummy_out_read -> fifo_dummy:avalonmm_read_slave_read
	signal mm_interconnect_1_switches_s1_readdata                                : std_logic_vector(31 downto 0);  -- switches:readdata -> mm_interconnect_1:switches_s1_readdata
	signal mm_interconnect_1_switches_s1_address                                 : std_logic_vector(1 downto 0);   -- mm_interconnect_1:switches_s1_address -> switches:address
	signal mm_interconnect_1_sdram_s1_chipselect                                 : std_logic;                      -- mm_interconnect_1:sdram_s1_chipselect -> sdram:az_cs
	signal mm_interconnect_1_sdram_s1_readdata                                   : std_logic_vector(15 downto 0);  -- sdram:za_data -> mm_interconnect_1:sdram_s1_readdata
	signal mm_interconnect_1_sdram_s1_waitrequest                                : std_logic;                      -- sdram:za_waitrequest -> mm_interconnect_1:sdram_s1_waitrequest
	signal mm_interconnect_1_sdram_s1_address                                    : std_logic_vector(24 downto 0);  -- mm_interconnect_1:sdram_s1_address -> sdram:az_addr
	signal mm_interconnect_1_sdram_s1_read                                       : std_logic;                      -- mm_interconnect_1:sdram_s1_read -> mm_interconnect_1_sdram_s1_read:in
	signal mm_interconnect_1_sdram_s1_byteenable                                 : std_logic_vector(1 downto 0);   -- mm_interconnect_1:sdram_s1_byteenable -> mm_interconnect_1_sdram_s1_byteenable:in
	signal mm_interconnect_1_sdram_s1_readdatavalid                              : std_logic;                      -- sdram:za_valid -> mm_interconnect_1:sdram_s1_readdatavalid
	signal mm_interconnect_1_sdram_s1_write                                      : std_logic;                      -- mm_interconnect_1:sdram_s1_write -> mm_interconnect_1_sdram_s1_write:in
	signal mm_interconnect_1_sdram_s1_writedata                                  : std_logic_vector(15 downto 0);  -- mm_interconnect_1:sdram_s1_writedata -> sdram:az_data
	signal mm_interconnect_1_adc_fifo_mem_out_readdata                           : std_logic_vector(31 downto 0);  -- adc_fifo_mem:avalonmm_read_slave_readdata -> mm_interconnect_1:adc_fifo_mem_out_readdata
	signal mm_interconnect_1_adc_fifo_mem_out_waitrequest                        : std_logic;                      -- adc_fifo_mem:avalonmm_read_slave_waitrequest -> mm_interconnect_1:adc_fifo_mem_out_waitrequest
	signal mm_interconnect_1_adc_fifo_mem_out_address                            : std_logic_vector(0 downto 0);   -- mm_interconnect_1:adc_fifo_mem_out_address -> adc_fifo_mem:avalonmm_read_slave_address
	signal mm_interconnect_1_adc_fifo_mem_out_read                               : std_logic;                      -- mm_interconnect_1:adc_fifo_mem_out_read -> adc_fifo_mem:avalonmm_read_slave_read
	signal mm_interconnect_1_nmr_parameters_adc_val_sub_s1_chipselect            : std_logic;                      -- mm_interconnect_1:nmr_parameters_adc_val_sub_s1_chipselect -> nmr_parameters:adc_val_sub_s1_chipselect
	signal mm_interconnect_1_nmr_parameters_adc_val_sub_s1_readdata              : std_logic_vector(31 downto 0);  -- nmr_parameters:adc_val_sub_s1_readdata -> mm_interconnect_1:nmr_parameters_adc_val_sub_s1_readdata
	signal mm_interconnect_1_nmr_parameters_adc_val_sub_s1_address               : std_logic_vector(1 downto 0);   -- mm_interconnect_1:nmr_parameters_adc_val_sub_s1_address -> nmr_parameters:adc_val_sub_s1_address
	signal mm_interconnect_1_nmr_parameters_adc_val_sub_s1_write                 : std_logic;                      -- mm_interconnect_1:nmr_parameters_adc_val_sub_s1_write -> mm_interconnect_1_nmr_parameters_adc_val_sub_s1_write:in
	signal mm_interconnect_1_nmr_parameters_adc_val_sub_s1_writedata             : std_logic_vector(31 downto 0);  -- mm_interconnect_1:nmr_parameters_adc_val_sub_s1_writedata -> nmr_parameters:adc_val_sub_s1_writedata
	signal mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect              : std_logic;                      -- mm_interconnect_1:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	signal mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata                : std_logic_vector(31 downto 0);  -- jtag_uart:av_readdata -> mm_interconnect_1:jtag_uart_avalon_jtag_slave_readdata
	signal mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest             : std_logic;                      -- jtag_uart:av_waitrequest -> mm_interconnect_1:jtag_uart_avalon_jtag_slave_waitrequest
	signal mm_interconnect_1_jtag_uart_avalon_jtag_slave_address                 : std_logic_vector(0 downto 0);   -- mm_interconnect_1:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	signal mm_interconnect_1_jtag_uart_avalon_jtag_slave_read                    : std_logic;                      -- mm_interconnect_1:jtag_uart_avalon_jtag_slave_read -> mm_interconnect_1_jtag_uart_avalon_jtag_slave_read:in
	signal mm_interconnect_1_jtag_uart_avalon_jtag_slave_write                   : std_logic;                      -- mm_interconnect_1:jtag_uart_avalon_jtag_slave_write -> mm_interconnect_1_jtag_uart_avalon_jtag_slave_write:in
	signal mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata               : std_logic_vector(31 downto 0);  -- mm_interconnect_1:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	signal mm_interconnect_1_dconv_fir_avalon_mm_slave_readdata                  : std_logic_vector(15 downto 0);  -- dconv_fir:coeff_out_data -> mm_interconnect_1:dconv_fir_avalon_mm_slave_readdata
	signal mm_interconnect_1_dconv_fir_avalon_mm_slave_address                   : std_logic_vector(5 downto 0);   -- mm_interconnect_1:dconv_fir_avalon_mm_slave_address -> dconv_fir:coeff_in_address
	signal mm_interconnect_1_dconv_fir_avalon_mm_slave_read                      : std_logic;                      -- mm_interconnect_1:dconv_fir_avalon_mm_slave_read -> dconv_fir:coeff_in_read
	signal mm_interconnect_1_dconv_fir_avalon_mm_slave_readdatavalid             : std_logic;                      -- dconv_fir:coeff_out_valid -> mm_interconnect_1:dconv_fir_avalon_mm_slave_readdatavalid
	signal mm_interconnect_1_dconv_fir_avalon_mm_slave_write                     : std_logic;                      -- mm_interconnect_1:dconv_fir_avalon_mm_slave_write -> dconv_fir:coeff_in_we
	signal mm_interconnect_1_dconv_fir_avalon_mm_slave_writedata                 : std_logic_vector(15 downto 0);  -- mm_interconnect_1:dconv_fir_avalon_mm_slave_writedata -> dconv_fir:coeff_in_data
	signal mm_interconnect_1_dconv_fir_q_avalon_mm_slave_readdata                : std_logic_vector(15 downto 0);  -- dconv_fir_q:coeff_out_data -> mm_interconnect_1:dconv_fir_q_avalon_mm_slave_readdata
	signal mm_interconnect_1_dconv_fir_q_avalon_mm_slave_address                 : std_logic_vector(5 downto 0);   -- mm_interconnect_1:dconv_fir_q_avalon_mm_slave_address -> dconv_fir_q:coeff_in_address
	signal mm_interconnect_1_dconv_fir_q_avalon_mm_slave_read                    : std_logic;                      -- mm_interconnect_1:dconv_fir_q_avalon_mm_slave_read -> dconv_fir_q:coeff_in_read
	signal mm_interconnect_1_dconv_fir_q_avalon_mm_slave_readdatavalid           : std_logic;                      -- dconv_fir_q:coeff_out_valid -> mm_interconnect_1:dconv_fir_q_avalon_mm_slave_readdatavalid
	signal mm_interconnect_1_dconv_fir_q_avalon_mm_slave_write                   : std_logic;                      -- mm_interconnect_1:dconv_fir_q_avalon_mm_slave_write -> dconv_fir_q:coeff_in_we
	signal mm_interconnect_1_dconv_fir_q_avalon_mm_slave_writedata               : std_logic_vector(15 downto 0);  -- mm_interconnect_1:dconv_fir_q_avalon_mm_slave_writedata -> dconv_fir_q:coeff_in_data
	signal mm_interconnect_1_alt_vip_vfr_vga_avalon_slave_readdata               : std_logic_vector(31 downto 0);  -- alt_vip_vfr_vga:slave_readdata -> mm_interconnect_1:alt_vip_vfr_vga_avalon_slave_readdata
	signal mm_interconnect_1_alt_vip_vfr_vga_avalon_slave_address                : std_logic_vector(4 downto 0);   -- mm_interconnect_1:alt_vip_vfr_vga_avalon_slave_address -> alt_vip_vfr_vga:slave_address
	signal mm_interconnect_1_alt_vip_vfr_vga_avalon_slave_read                   : std_logic;                      -- mm_interconnect_1:alt_vip_vfr_vga_avalon_slave_read -> alt_vip_vfr_vga:slave_read
	signal mm_interconnect_1_alt_vip_vfr_vga_avalon_slave_write                  : std_logic;                      -- mm_interconnect_1:alt_vip_vfr_vga_avalon_slave_write -> alt_vip_vfr_vga:slave_write
	signal mm_interconnect_1_alt_vip_vfr_vga_avalon_slave_writedata              : std_logic_vector(31 downto 0);  -- mm_interconnect_1:alt_vip_vfr_vga_avalon_slave_writedata -> alt_vip_vfr_vga:slave_writedata
	signal mm_interconnect_1_sysid_qsys_control_slave_readdata                   : std_logic_vector(31 downto 0);  -- sysid_qsys:readdata -> mm_interconnect_1:sysid_qsys_control_slave_readdata
	signal mm_interconnect_1_sysid_qsys_control_slave_address                    : std_logic_vector(0 downto 0);   -- mm_interconnect_1:sysid_qsys_control_slave_address -> sysid_qsys:address
	signal mm_interconnect_1_i2c_int_csr_readdata                                : std_logic_vector(31 downto 0);  -- i2c_int:readdata -> mm_interconnect_1:i2c_int_csr_readdata
	signal mm_interconnect_1_i2c_int_csr_address                                 : std_logic_vector(3 downto 0);   -- mm_interconnect_1:i2c_int_csr_address -> i2c_int:addr
	signal mm_interconnect_1_i2c_int_csr_read                                    : std_logic;                      -- mm_interconnect_1:i2c_int_csr_read -> i2c_int:read
	signal mm_interconnect_1_i2c_int_csr_write                                   : std_logic;                      -- mm_interconnect_1:i2c_int_csr_write -> i2c_int:write
	signal mm_interconnect_1_i2c_int_csr_writedata                               : std_logic_vector(31 downto 0);  -- mm_interconnect_1:i2c_int_csr_writedata -> i2c_int:writedata
	signal mm_interconnect_1_i2c_ext_csr_readdata                                : std_logic_vector(31 downto 0);  -- i2c_ext:readdata -> mm_interconnect_1:i2c_ext_csr_readdata
	signal mm_interconnect_1_i2c_ext_csr_address                                 : std_logic_vector(3 downto 0);   -- mm_interconnect_1:i2c_ext_csr_address -> i2c_ext:addr
	signal mm_interconnect_1_i2c_ext_csr_read                                    : std_logic;                      -- mm_interconnect_1:i2c_ext_csr_read -> i2c_ext:read
	signal mm_interconnect_1_i2c_ext_csr_write                                   : std_logic;                      -- mm_interconnect_1:i2c_ext_csr_write -> i2c_ext:write
	signal mm_interconnect_1_i2c_ext_csr_writedata                               : std_logic_vector(31 downto 0);  -- mm_interconnect_1:i2c_ext_csr_writedata -> i2c_ext:writedata
	signal mm_interconnect_1_nmr_parameters_delay_nosig_s1_chipselect            : std_logic;                      -- mm_interconnect_1:nmr_parameters_delay_nosig_s1_chipselect -> nmr_parameters:delay_nosig_s1_chipselect
	signal mm_interconnect_1_nmr_parameters_delay_nosig_s1_readdata              : std_logic_vector(31 downto 0);  -- nmr_parameters:delay_nosig_s1_readdata -> mm_interconnect_1:nmr_parameters_delay_nosig_s1_readdata
	signal mm_interconnect_1_nmr_parameters_delay_nosig_s1_address               : std_logic_vector(1 downto 0);   -- mm_interconnect_1:nmr_parameters_delay_nosig_s1_address -> nmr_parameters:delay_nosig_s1_address
	signal mm_interconnect_1_nmr_parameters_delay_nosig_s1_write                 : std_logic;                      -- mm_interconnect_1:nmr_parameters_delay_nosig_s1_write -> mm_interconnect_1_nmr_parameters_delay_nosig_s1_write:in
	signal mm_interconnect_1_nmr_parameters_delay_nosig_s1_writedata             : std_logic_vector(31 downto 0);  -- mm_interconnect_1:nmr_parameters_delay_nosig_s1_writedata -> nmr_parameters:delay_nosig_s1_writedata
	signal mm_interconnect_1_nmr_parameters_delay_sig_s1_chipselect              : std_logic;                      -- mm_interconnect_1:nmr_parameters_delay_sig_s1_chipselect -> nmr_parameters:delay_sig_s1_chipselect
	signal mm_interconnect_1_nmr_parameters_delay_sig_s1_readdata                : std_logic_vector(31 downto 0);  -- nmr_parameters:delay_sig_s1_readdata -> mm_interconnect_1:nmr_parameters_delay_sig_s1_readdata
	signal mm_interconnect_1_nmr_parameters_delay_sig_s1_address                 : std_logic_vector(1 downto 0);   -- mm_interconnect_1:nmr_parameters_delay_sig_s1_address -> nmr_parameters:delay_sig_s1_address
	signal mm_interconnect_1_nmr_parameters_delay_sig_s1_write                   : std_logic;                      -- mm_interconnect_1:nmr_parameters_delay_sig_s1_write -> mm_interconnect_1_nmr_parameters_delay_sig_s1_write:in
	signal mm_interconnect_1_nmr_parameters_delay_sig_s1_writedata               : std_logic_vector(31 downto 0);  -- mm_interconnect_1:nmr_parameters_delay_sig_s1_writedata -> nmr_parameters:delay_sig_s1_writedata
	signal mm_interconnect_1_nmr_parameters_delay_t1_s1_chipselect               : std_logic;                      -- mm_interconnect_1:nmr_parameters_delay_t1_s1_chipselect -> nmr_parameters:delay_t1_s1_chipselect
	signal mm_interconnect_1_nmr_parameters_delay_t1_s1_readdata                 : std_logic_vector(31 downto 0);  -- nmr_parameters:delay_t1_s1_readdata -> mm_interconnect_1:nmr_parameters_delay_t1_s1_readdata
	signal mm_interconnect_1_nmr_parameters_delay_t1_s1_address                  : std_logic_vector(1 downto 0);   -- mm_interconnect_1:nmr_parameters_delay_t1_s1_address -> nmr_parameters:delay_t1_s1_address
	signal mm_interconnect_1_nmr_parameters_delay_t1_s1_write                    : std_logic;                      -- mm_interconnect_1:nmr_parameters_delay_t1_s1_write -> mm_interconnect_1_nmr_parameters_delay_t1_s1_write:in
	signal mm_interconnect_1_nmr_parameters_delay_t1_s1_writedata                : std_logic_vector(31 downto 0);  -- mm_interconnect_1:nmr_parameters_delay_t1_s1_writedata -> nmr_parameters:delay_t1_s1_writedata
	signal mm_interconnect_1_nmr_parameters_echoes_per_scan_s1_chipselect        : std_logic;                      -- mm_interconnect_1:nmr_parameters_echoes_per_scan_s1_chipselect -> nmr_parameters:echoes_per_scan_s1_chipselect
	signal mm_interconnect_1_nmr_parameters_echoes_per_scan_s1_readdata          : std_logic_vector(31 downto 0);  -- nmr_parameters:echoes_per_scan_s1_readdata -> mm_interconnect_1:nmr_parameters_echoes_per_scan_s1_readdata
	signal mm_interconnect_1_nmr_parameters_echoes_per_scan_s1_address           : std_logic_vector(1 downto 0);   -- mm_interconnect_1:nmr_parameters_echoes_per_scan_s1_address -> nmr_parameters:echoes_per_scan_s1_address
	signal mm_interconnect_1_nmr_parameters_echoes_per_scan_s1_write             : std_logic;                      -- mm_interconnect_1:nmr_parameters_echoes_per_scan_s1_write -> mm_interconnect_1_nmr_parameters_echoes_per_scan_s1_write:in
	signal mm_interconnect_1_nmr_parameters_echoes_per_scan_s1_writedata         : std_logic_vector(31 downto 0);  -- mm_interconnect_1:nmr_parameters_echoes_per_scan_s1_writedata -> nmr_parameters:echoes_per_scan_s1_writedata
	signal mm_interconnect_1_adc_fifo_mem_in_csr_readdata                        : std_logic_vector(31 downto 0);  -- adc_fifo_mem:wrclk_control_slave_readdata -> mm_interconnect_1:adc_fifo_mem_in_csr_readdata
	signal mm_interconnect_1_adc_fifo_mem_in_csr_address                         : std_logic_vector(2 downto 0);   -- mm_interconnect_1:adc_fifo_mem_in_csr_address -> adc_fifo_mem:wrclk_control_slave_address
	signal mm_interconnect_1_adc_fifo_mem_in_csr_read                            : std_logic;                      -- mm_interconnect_1:adc_fifo_mem_in_csr_read -> adc_fifo_mem:wrclk_control_slave_read
	signal mm_interconnect_1_adc_fifo_mem_in_csr_write                           : std_logic;                      -- mm_interconnect_1:adc_fifo_mem_in_csr_write -> adc_fifo_mem:wrclk_control_slave_write
	signal mm_interconnect_1_adc_fifo_mem_in_csr_writedata                       : std_logic_vector(31 downto 0);  -- mm_interconnect_1:adc_fifo_mem_in_csr_writedata -> adc_fifo_mem:wrclk_control_slave_writedata
	signal mm_interconnect_1_dconv_fifo_mem_in_csr_readdata                      : std_logic_vector(31 downto 0);  -- dconv_fifo_mem:wrclk_control_slave_readdata -> mm_interconnect_1:dconv_fifo_mem_in_csr_readdata
	signal mm_interconnect_1_dconv_fifo_mem_in_csr_address                       : std_logic_vector(2 downto 0);   -- mm_interconnect_1:dconv_fifo_mem_in_csr_address -> dconv_fifo_mem:wrclk_control_slave_address
	signal mm_interconnect_1_dconv_fifo_mem_in_csr_read                          : std_logic;                      -- mm_interconnect_1:dconv_fifo_mem_in_csr_read -> dconv_fifo_mem:wrclk_control_slave_read
	signal mm_interconnect_1_dconv_fifo_mem_in_csr_write                         : std_logic;                      -- mm_interconnect_1:dconv_fifo_mem_in_csr_write -> dconv_fifo_mem:wrclk_control_slave_write
	signal mm_interconnect_1_dconv_fifo_mem_in_csr_writedata                     : std_logic_vector(31 downto 0);  -- mm_interconnect_1:dconv_fifo_mem_in_csr_writedata -> dconv_fifo_mem:wrclk_control_slave_writedata
	signal mm_interconnect_1_dconv_fifo_mem_q_in_csr_readdata                    : std_logic_vector(31 downto 0);  -- dconv_fifo_mem_q:wrclk_control_slave_readdata -> mm_interconnect_1:dconv_fifo_mem_q_in_csr_readdata
	signal mm_interconnect_1_dconv_fifo_mem_q_in_csr_address                     : std_logic_vector(2 downto 0);   -- mm_interconnect_1:dconv_fifo_mem_q_in_csr_address -> dconv_fifo_mem_q:wrclk_control_slave_address
	signal mm_interconnect_1_dconv_fifo_mem_q_in_csr_read                        : std_logic;                      -- mm_interconnect_1:dconv_fifo_mem_q_in_csr_read -> dconv_fifo_mem_q:wrclk_control_slave_read
	signal mm_interconnect_1_dconv_fifo_mem_q_in_csr_write                       : std_logic;                      -- mm_interconnect_1:dconv_fifo_mem_q_in_csr_write -> dconv_fifo_mem_q:wrclk_control_slave_write
	signal mm_interconnect_1_dconv_fifo_mem_q_in_csr_writedata                   : std_logic_vector(31 downto 0);  -- mm_interconnect_1:dconv_fifo_mem_q_in_csr_writedata -> dconv_fifo_mem_q:wrclk_control_slave_writedata
	signal mm_interconnect_1_nmr_parameters_init_delay_s1_chipselect             : std_logic;                      -- mm_interconnect_1:nmr_parameters_init_delay_s1_chipselect -> nmr_parameters:init_delay_s1_chipselect
	signal mm_interconnect_1_nmr_parameters_init_delay_s1_readdata               : std_logic_vector(31 downto 0);  -- nmr_parameters:init_delay_s1_readdata -> mm_interconnect_1:nmr_parameters_init_delay_s1_readdata
	signal mm_interconnect_1_nmr_parameters_init_delay_s1_address                : std_logic_vector(1 downto 0);   -- mm_interconnect_1:nmr_parameters_init_delay_s1_address -> nmr_parameters:init_delay_s1_address
	signal mm_interconnect_1_nmr_parameters_init_delay_s1_write                  : std_logic;                      -- mm_interconnect_1:nmr_parameters_init_delay_s1_write -> mm_interconnect_1_nmr_parameters_init_delay_s1_write:in
	signal mm_interconnect_1_nmr_parameters_init_delay_s1_writedata              : std_logic_vector(31 downto 0);  -- mm_interconnect_1:nmr_parameters_init_delay_s1_writedata -> nmr_parameters:init_delay_s1_writedata
	signal mm_interconnect_1_nmr_sys_pll_reconfig_mgmt_avalon_slave_readdata     : std_logic_vector(31 downto 0);  -- nmr_sys_pll_reconfig:mgmt_readdata -> mm_interconnect_1:nmr_sys_pll_reconfig_mgmt_avalon_slave_readdata
	signal mm_interconnect_1_nmr_sys_pll_reconfig_mgmt_avalon_slave_waitrequest  : std_logic;                      -- nmr_sys_pll_reconfig:mgmt_waitrequest -> mm_interconnect_1:nmr_sys_pll_reconfig_mgmt_avalon_slave_waitrequest
	signal mm_interconnect_1_nmr_sys_pll_reconfig_mgmt_avalon_slave_address      : std_logic_vector(5 downto 0);   -- mm_interconnect_1:nmr_sys_pll_reconfig_mgmt_avalon_slave_address -> nmr_sys_pll_reconfig:mgmt_address
	signal mm_interconnect_1_nmr_sys_pll_reconfig_mgmt_avalon_slave_read         : std_logic;                      -- mm_interconnect_1:nmr_sys_pll_reconfig_mgmt_avalon_slave_read -> nmr_sys_pll_reconfig:mgmt_read
	signal mm_interconnect_1_nmr_sys_pll_reconfig_mgmt_avalon_slave_write        : std_logic;                      -- mm_interconnect_1:nmr_sys_pll_reconfig_mgmt_avalon_slave_write -> nmr_sys_pll_reconfig:mgmt_write
	signal mm_interconnect_1_nmr_sys_pll_reconfig_mgmt_avalon_slave_writedata    : std_logic_vector(31 downto 0);  -- mm_interconnect_1:nmr_sys_pll_reconfig_mgmt_avalon_slave_writedata -> nmr_sys_pll_reconfig:mgmt_writedata
	signal mm_interconnect_1_analyzer_pll_reconfig_mgmt_avalon_slave_readdata    : std_logic_vector(31 downto 0);  -- analyzer_pll_reconfig:mgmt_readdata -> mm_interconnect_1:analyzer_pll_reconfig_mgmt_avalon_slave_readdata
	signal mm_interconnect_1_analyzer_pll_reconfig_mgmt_avalon_slave_waitrequest : std_logic;                      -- analyzer_pll_reconfig:mgmt_waitrequest -> mm_interconnect_1:analyzer_pll_reconfig_mgmt_avalon_slave_waitrequest
	signal mm_interconnect_1_analyzer_pll_reconfig_mgmt_avalon_slave_address     : std_logic_vector(5 downto 0);   -- mm_interconnect_1:analyzer_pll_reconfig_mgmt_avalon_slave_address -> analyzer_pll_reconfig:mgmt_address
	signal mm_interconnect_1_analyzer_pll_reconfig_mgmt_avalon_slave_read        : std_logic;                      -- mm_interconnect_1:analyzer_pll_reconfig_mgmt_avalon_slave_read -> analyzer_pll_reconfig:mgmt_read
	signal mm_interconnect_1_analyzer_pll_reconfig_mgmt_avalon_slave_write       : std_logic;                      -- mm_interconnect_1:analyzer_pll_reconfig_mgmt_avalon_slave_write -> analyzer_pll_reconfig:mgmt_write
	signal mm_interconnect_1_analyzer_pll_reconfig_mgmt_avalon_slave_writedata   : std_logic_vector(31 downto 0);  -- mm_interconnect_1:analyzer_pll_reconfig_mgmt_avalon_slave_writedata -> analyzer_pll_reconfig:mgmt_writedata
	signal mm_interconnect_1_dconv_fifo_mem_out_readdata                         : std_logic_vector(31 downto 0);  -- dconv_fifo_mem:avalonmm_read_slave_readdata -> mm_interconnect_1:dconv_fifo_mem_out_readdata
	signal mm_interconnect_1_dconv_fifo_mem_out_waitrequest                      : std_logic;                      -- dconv_fifo_mem:avalonmm_read_slave_waitrequest -> mm_interconnect_1:dconv_fifo_mem_out_waitrequest
	signal mm_interconnect_1_dconv_fifo_mem_out_address                          : std_logic_vector(0 downto 0);   -- mm_interconnect_1:dconv_fifo_mem_out_address -> dconv_fifo_mem:avalonmm_read_slave_address
	signal mm_interconnect_1_dconv_fifo_mem_out_read                             : std_logic;                      -- mm_interconnect_1:dconv_fifo_mem_out_read -> dconv_fifo_mem:avalonmm_read_slave_read
	signal mm_interconnect_1_dconv_fifo_mem_q_out_readdata                       : std_logic_vector(31 downto 0);  -- dconv_fifo_mem_q:avalonmm_read_slave_readdata -> mm_interconnect_1:dconv_fifo_mem_q_out_readdata
	signal mm_interconnect_1_dconv_fifo_mem_q_out_waitrequest                    : std_logic;                      -- dconv_fifo_mem_q:avalonmm_read_slave_waitrequest -> mm_interconnect_1:dconv_fifo_mem_q_out_waitrequest
	signal mm_interconnect_1_dconv_fifo_mem_q_out_address                        : std_logic_vector(0 downto 0);   -- mm_interconnect_1:dconv_fifo_mem_q_out_address -> dconv_fifo_mem_q:avalonmm_read_slave_address
	signal mm_interconnect_1_dconv_fifo_mem_q_out_read                           : std_logic;                      -- mm_interconnect_1:dconv_fifo_mem_q_out_read -> dconv_fifo_mem_q:avalonmm_read_slave_read
	signal mm_interconnect_1_nmr_parameters_pulse_180deg_s1_chipselect           : std_logic;                      -- mm_interconnect_1:nmr_parameters_pulse_180deg_s1_chipselect -> nmr_parameters:pulse_180deg_s1_chipselect
	signal mm_interconnect_1_nmr_parameters_pulse_180deg_s1_readdata             : std_logic_vector(31 downto 0);  -- nmr_parameters:pulse_180deg_s1_readdata -> mm_interconnect_1:nmr_parameters_pulse_180deg_s1_readdata
	signal mm_interconnect_1_nmr_parameters_pulse_180deg_s1_address              : std_logic_vector(1 downto 0);   -- mm_interconnect_1:nmr_parameters_pulse_180deg_s1_address -> nmr_parameters:pulse_180deg_s1_address
	signal mm_interconnect_1_nmr_parameters_pulse_180deg_s1_write                : std_logic;                      -- mm_interconnect_1:nmr_parameters_pulse_180deg_s1_write -> mm_interconnect_1_nmr_parameters_pulse_180deg_s1_write:in
	signal mm_interconnect_1_nmr_parameters_pulse_180deg_s1_writedata            : std_logic_vector(31 downto 0);  -- mm_interconnect_1:nmr_parameters_pulse_180deg_s1_writedata -> nmr_parameters:pulse_180deg_s1_writedata
	signal mm_interconnect_1_nmr_parameters_pulse_90deg_s1_chipselect            : std_logic;                      -- mm_interconnect_1:nmr_parameters_pulse_90deg_s1_chipselect -> nmr_parameters:pulse_90deg_s1_chipselect
	signal mm_interconnect_1_nmr_parameters_pulse_90deg_s1_readdata              : std_logic_vector(31 downto 0);  -- nmr_parameters:pulse_90deg_s1_readdata -> mm_interconnect_1:nmr_parameters_pulse_90deg_s1_readdata
	signal mm_interconnect_1_nmr_parameters_pulse_90deg_s1_address               : std_logic_vector(1 downto 0);   -- mm_interconnect_1:nmr_parameters_pulse_90deg_s1_address -> nmr_parameters:pulse_90deg_s1_address
	signal mm_interconnect_1_nmr_parameters_pulse_90deg_s1_write                 : std_logic;                      -- mm_interconnect_1:nmr_parameters_pulse_90deg_s1_write -> mm_interconnect_1_nmr_parameters_pulse_90deg_s1_write:in
	signal mm_interconnect_1_nmr_parameters_pulse_90deg_s1_writedata             : std_logic_vector(31 downto 0);  -- mm_interconnect_1:nmr_parameters_pulse_90deg_s1_writedata -> nmr_parameters:pulse_90deg_s1_writedata
	signal mm_interconnect_1_nmr_parameters_pulse_t1_s1_chipselect               : std_logic;                      -- mm_interconnect_1:nmr_parameters_pulse_t1_s1_chipselect -> nmr_parameters:pulse_t1_s1_chipselect
	signal mm_interconnect_1_nmr_parameters_pulse_t1_s1_readdata                 : std_logic_vector(31 downto 0);  -- nmr_parameters:pulse_t1_s1_readdata -> mm_interconnect_1:nmr_parameters_pulse_t1_s1_readdata
	signal mm_interconnect_1_nmr_parameters_pulse_t1_s1_address                  : std_logic_vector(1 downto 0);   -- mm_interconnect_1:nmr_parameters_pulse_t1_s1_address -> nmr_parameters:pulse_t1_s1_address
	signal mm_interconnect_1_nmr_parameters_pulse_t1_s1_write                    : std_logic;                      -- mm_interconnect_1:nmr_parameters_pulse_t1_s1_write -> mm_interconnect_1_nmr_parameters_pulse_t1_s1_write:in
	signal mm_interconnect_1_nmr_parameters_pulse_t1_s1_writedata                : std_logic_vector(31 downto 0);  -- mm_interconnect_1:nmr_parameters_pulse_t1_s1_writedata -> nmr_parameters:pulse_t1_s1_writedata
	signal mm_interconnect_1_nmr_parameters_rx_delay_s1_chipselect               : std_logic;                      -- mm_interconnect_1:nmr_parameters_rx_delay_s1_chipselect -> nmr_parameters:rx_delay_s1_chipselect
	signal mm_interconnect_1_nmr_parameters_rx_delay_s1_readdata                 : std_logic_vector(31 downto 0);  -- nmr_parameters:rx_delay_s1_readdata -> mm_interconnect_1:nmr_parameters_rx_delay_s1_readdata
	signal mm_interconnect_1_nmr_parameters_rx_delay_s1_address                  : std_logic_vector(1 downto 0);   -- mm_interconnect_1:nmr_parameters_rx_delay_s1_address -> nmr_parameters:rx_delay_s1_address
	signal mm_interconnect_1_nmr_parameters_rx_delay_s1_write                    : std_logic;                      -- mm_interconnect_1:nmr_parameters_rx_delay_s1_write -> mm_interconnect_1_nmr_parameters_rx_delay_s1_write:in
	signal mm_interconnect_1_nmr_parameters_rx_delay_s1_writedata                : std_logic_vector(31 downto 0);  -- mm_interconnect_1:nmr_parameters_rx_delay_s1_writedata -> nmr_parameters:rx_delay_s1_writedata
	signal mm_interconnect_1_ctrl_out_s1_chipselect                              : std_logic;                      -- mm_interconnect_1:ctrl_out_s1_chipselect -> ctrl_out:chipselect
	signal mm_interconnect_1_ctrl_out_s1_readdata                                : std_logic_vector(31 downto 0);  -- ctrl_out:readdata -> mm_interconnect_1:ctrl_out_s1_readdata
	signal mm_interconnect_1_ctrl_out_s1_address                                 : std_logic_vector(1 downto 0);   -- mm_interconnect_1:ctrl_out_s1_address -> ctrl_out:address
	signal mm_interconnect_1_ctrl_out_s1_write                                   : std_logic;                      -- mm_interconnect_1:ctrl_out_s1_write -> mm_interconnect_1_ctrl_out_s1_write:in
	signal mm_interconnect_1_ctrl_out_s1_writedata                               : std_logic_vector(31 downto 0);  -- mm_interconnect_1:ctrl_out_s1_writedata -> ctrl_out:writedata
	signal mm_interconnect_1_ctrl_in_s1_readdata                                 : std_logic_vector(31 downto 0);  -- ctrl_in:readdata -> mm_interconnect_1:ctrl_in_s1_readdata
	signal mm_interconnect_1_ctrl_in_s1_address                                  : std_logic_vector(1 downto 0);   -- mm_interconnect_1:ctrl_in_s1_address -> ctrl_in:address
	signal mm_interconnect_1_aux_cnt_out_s1_chipselect                           : std_logic;                      -- mm_interconnect_1:aux_cnt_out_s1_chipselect -> aux_cnt_out:chipselect
	signal mm_interconnect_1_aux_cnt_out_s1_readdata                             : std_logic_vector(31 downto 0);  -- aux_cnt_out:readdata -> mm_interconnect_1:aux_cnt_out_s1_readdata
	signal mm_interconnect_1_aux_cnt_out_s1_address                              : std_logic_vector(1 downto 0);   -- mm_interconnect_1:aux_cnt_out_s1_address -> aux_cnt_out:address
	signal mm_interconnect_1_aux_cnt_out_s1_write                                : std_logic;                      -- mm_interconnect_1:aux_cnt_out_s1_write -> mm_interconnect_1_aux_cnt_out_s1_write:in
	signal mm_interconnect_1_aux_cnt_out_s1_writedata                            : std_logic_vector(31 downto 0);  -- mm_interconnect_1:aux_cnt_out_s1_writedata -> aux_cnt_out:writedata
	signal mm_interconnect_1_nmr_parameters_samples_per_echo_s1_chipselect       : std_logic;                      -- mm_interconnect_1:nmr_parameters_samples_per_echo_s1_chipselect -> nmr_parameters:samples_per_echo_s1_chipselect
	signal mm_interconnect_1_nmr_parameters_samples_per_echo_s1_readdata         : std_logic_vector(31 downto 0);  -- nmr_parameters:samples_per_echo_s1_readdata -> mm_interconnect_1:nmr_parameters_samples_per_echo_s1_readdata
	signal mm_interconnect_1_nmr_parameters_samples_per_echo_s1_address          : std_logic_vector(1 downto 0);   -- mm_interconnect_1:nmr_parameters_samples_per_echo_s1_address -> nmr_parameters:samples_per_echo_s1_address
	signal mm_interconnect_1_nmr_parameters_samples_per_echo_s1_write            : std_logic;                      -- mm_interconnect_1:nmr_parameters_samples_per_echo_s1_write -> mm_interconnect_1_nmr_parameters_samples_per_echo_s1_write:in
	signal mm_interconnect_1_nmr_parameters_samples_per_echo_s1_writedata        : std_logic_vector(31 downto 0);  -- mm_interconnect_1:nmr_parameters_samples_per_echo_s1_writedata -> nmr_parameters:samples_per_echo_s1_writedata
	signal mm_interconnect_1_dac_grad_spi_control_port_chipselect                : std_logic;                      -- mm_interconnect_1:dac_grad_spi_control_port_chipselect -> dac_grad:spi_select
	signal mm_interconnect_1_dac_grad_spi_control_port_readdata                  : std_logic_vector(31 downto 0);  -- dac_grad:data_to_cpu -> mm_interconnect_1:dac_grad_spi_control_port_readdata
	signal mm_interconnect_1_dac_grad_spi_control_port_address                   : std_logic_vector(2 downto 0);   -- mm_interconnect_1:dac_grad_spi_control_port_address -> dac_grad:mem_addr
	signal mm_interconnect_1_dac_grad_spi_control_port_read                      : std_logic;                      -- mm_interconnect_1:dac_grad_spi_control_port_read -> mm_interconnect_1_dac_grad_spi_control_port_read:in
	signal mm_interconnect_1_dac_grad_spi_control_port_write                     : std_logic;                      -- mm_interconnect_1:dac_grad_spi_control_port_write -> mm_interconnect_1_dac_grad_spi_control_port_write:in
	signal mm_interconnect_1_dac_grad_spi_control_port_writedata                 : std_logic_vector(31 downto 0);  -- mm_interconnect_1:dac_grad_spi_control_port_writedata -> dac_grad:data_from_cpu
	signal mm_interconnect_1_spi_mtch_ntwrk_spi_control_port_chipselect          : std_logic;                      -- mm_interconnect_1:spi_mtch_ntwrk_spi_control_port_chipselect -> spi_mtch_ntwrk:spi_select
	signal mm_interconnect_1_spi_mtch_ntwrk_spi_control_port_readdata            : std_logic_vector(31 downto 0);  -- spi_mtch_ntwrk:data_to_cpu -> mm_interconnect_1:spi_mtch_ntwrk_spi_control_port_readdata
	signal mm_interconnect_1_spi_mtch_ntwrk_spi_control_port_address             : std_logic_vector(2 downto 0);   -- mm_interconnect_1:spi_mtch_ntwrk_spi_control_port_address -> spi_mtch_ntwrk:mem_addr
	signal mm_interconnect_1_spi_mtch_ntwrk_spi_control_port_read                : std_logic;                      -- mm_interconnect_1:spi_mtch_ntwrk_spi_control_port_read -> mm_interconnect_1_spi_mtch_ntwrk_spi_control_port_read:in
	signal mm_interconnect_1_spi_mtch_ntwrk_spi_control_port_write               : std_logic;                      -- mm_interconnect_1:spi_mtch_ntwrk_spi_control_port_write -> mm_interconnect_1_spi_mtch_ntwrk_spi_control_port_write:in
	signal mm_interconnect_1_spi_mtch_ntwrk_spi_control_port_writedata           : std_logic_vector(31 downto 0);  -- mm_interconnect_1:spi_mtch_ntwrk_spi_control_port_writedata -> spi_mtch_ntwrk:data_from_cpu
	signal mm_interconnect_1_spi_afe_relays_spi_control_port_chipselect          : std_logic;                      -- mm_interconnect_1:spi_afe_relays_spi_control_port_chipselect -> spi_afe_relays:spi_select
	signal mm_interconnect_1_spi_afe_relays_spi_control_port_readdata            : std_logic_vector(31 downto 0);  -- spi_afe_relays:data_to_cpu -> mm_interconnect_1:spi_afe_relays_spi_control_port_readdata
	signal mm_interconnect_1_spi_afe_relays_spi_control_port_address             : std_logic_vector(2 downto 0);   -- mm_interconnect_1:spi_afe_relays_spi_control_port_address -> spi_afe_relays:mem_addr
	signal mm_interconnect_1_spi_afe_relays_spi_control_port_read                : std_logic;                      -- mm_interconnect_1:spi_afe_relays_spi_control_port_read -> mm_interconnect_1_spi_afe_relays_spi_control_port_read:in
	signal mm_interconnect_1_spi_afe_relays_spi_control_port_write               : std_logic;                      -- mm_interconnect_1:spi_afe_relays_spi_control_port_write -> mm_interconnect_1_spi_afe_relays_spi_control_port_write:in
	signal mm_interconnect_1_spi_afe_relays_spi_control_port_writedata           : std_logic_vector(31 downto 0);  -- mm_interconnect_1:spi_afe_relays_spi_control_port_writedata -> spi_afe_relays:data_from_cpu
	signal mm_interconnect_1_dma_fifo_control_port_slave_chipselect              : std_logic;                      -- mm_interconnect_1:dma_fifo_control_port_slave_chipselect -> dma_fifo:dma_ctl_chipselect
	signal mm_interconnect_1_dma_fifo_control_port_slave_readdata                : std_logic_vector(31 downto 0);  -- dma_fifo:dma_ctl_readdata -> mm_interconnect_1:dma_fifo_control_port_slave_readdata
	signal mm_interconnect_1_dma_fifo_control_port_slave_address                 : std_logic_vector(2 downto 0);   -- mm_interconnect_1:dma_fifo_control_port_slave_address -> dma_fifo:dma_ctl_address
	signal mm_interconnect_1_dma_fifo_control_port_slave_write                   : std_logic;                      -- mm_interconnect_1:dma_fifo_control_port_slave_write -> mm_interconnect_1_dma_fifo_control_port_slave_write:in
	signal mm_interconnect_1_dma_fifo_control_port_slave_writedata               : std_logic_vector(31 downto 0);  -- mm_interconnect_1:dma_fifo_control_port_slave_writedata -> dma_fifo:dma_ctl_writedata
	signal mm_interconnect_1_dma_dconvi_control_port_slave_chipselect            : std_logic;                      -- mm_interconnect_1:dma_dconvi_control_port_slave_chipselect -> dma_dconvi:dma_ctl_chipselect
	signal mm_interconnect_1_dma_dconvi_control_port_slave_readdata              : std_logic_vector(31 downto 0);  -- dma_dconvi:dma_ctl_readdata -> mm_interconnect_1:dma_dconvi_control_port_slave_readdata
	signal mm_interconnect_1_dma_dconvi_control_port_slave_address               : std_logic_vector(2 downto 0);   -- mm_interconnect_1:dma_dconvi_control_port_slave_address -> dma_dconvi:dma_ctl_address
	signal mm_interconnect_1_dma_dconvi_control_port_slave_write                 : std_logic;                      -- mm_interconnect_1:dma_dconvi_control_port_slave_write -> mm_interconnect_1_dma_dconvi_control_port_slave_write:in
	signal mm_interconnect_1_dma_dconvi_control_port_slave_writedata             : std_logic_vector(31 downto 0);  -- mm_interconnect_1:dma_dconvi_control_port_slave_writedata -> dma_dconvi:dma_ctl_writedata
	signal mm_interconnect_1_dma_dconvq_control_port_slave_chipselect            : std_logic;                      -- mm_interconnect_1:dma_dconvq_control_port_slave_chipselect -> dma_dconvq:dma_ctl_chipselect
	signal mm_interconnect_1_dma_dconvq_control_port_slave_readdata              : std_logic_vector(31 downto 0);  -- dma_dconvq:dma_ctl_readdata -> mm_interconnect_1:dma_dconvq_control_port_slave_readdata
	signal mm_interconnect_1_dma_dconvq_control_port_slave_address               : std_logic_vector(2 downto 0);   -- mm_interconnect_1:dma_dconvq_control_port_slave_address -> dma_dconvq:dma_ctl_address
	signal mm_interconnect_1_dma_dconvq_control_port_slave_write                 : std_logic;                      -- mm_interconnect_1:dma_dconvq_control_port_slave_write -> mm_interconnect_1_dma_dconvq_control_port_slave_write:in
	signal mm_interconnect_1_dma_dconvq_control_port_slave_writedata             : std_logic_vector(31 downto 0);  -- mm_interconnect_1:dma_dconvq_control_port_slave_writedata -> dma_dconvq:dma_ctl_writedata
	signal mm_interconnect_1_dma_dummy_control_port_slave_chipselect             : std_logic;                      -- mm_interconnect_1:dma_dummy_control_port_slave_chipselect -> dma_dummy:dma_ctl_chipselect
	signal mm_interconnect_1_dma_dummy_control_port_slave_readdata               : std_logic_vector(31 downto 0);  -- dma_dummy:dma_ctl_readdata -> mm_interconnect_1:dma_dummy_control_port_slave_readdata
	signal mm_interconnect_1_dma_dummy_control_port_slave_address                : std_logic_vector(2 downto 0);   -- mm_interconnect_1:dma_dummy_control_port_slave_address -> dma_dummy:dma_ctl_address
	signal mm_interconnect_1_dma_dummy_control_port_slave_write                  : std_logic;                      -- mm_interconnect_1:dma_dummy_control_port_slave_write -> mm_interconnect_1_dma_dummy_control_port_slave_write:in
	signal mm_interconnect_1_dma_dummy_control_port_slave_writedata              : std_logic_vector(31 downto 0);  -- mm_interconnect_1:dma_dummy_control_port_slave_writedata -> dma_dummy:dma_ctl_writedata
	signal irq_mapper_receiver0_irq                                              : std_logic;                      -- alt_vip_vfr_vga:slave_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                              : std_logic;                      -- jtag_uart:av_irq -> irq_mapper:receiver1_irq
	signal hps_0_f2h_irq0_irq                                                    : std_logic_vector(31 downto 0);  -- irq_mapper:sender_irq -> hps_0:f2h_irq_p0
	signal irq_mapper_001_receiver0_irq                                          : std_logic;                      -- i2c_int:intr -> irq_mapper_001:receiver0_irq
	signal irq_mapper_001_receiver1_irq                                          : std_logic;                      -- i2c_ext:intr -> irq_mapper_001:receiver1_irq
	signal irq_mapper_001_receiver2_irq                                          : std_logic;                      -- dac_grad:irq -> irq_mapper_001:receiver2_irq
	signal irq_mapper_001_receiver3_irq                                          : std_logic;                      -- dma_fifo:dma_ctl_irq -> irq_mapper_001:receiver3_irq
	signal irq_mapper_001_receiver4_irq                                          : std_logic;                      -- spi_mtch_ntwrk:irq -> irq_mapper_001:receiver4_irq
	signal irq_mapper_001_receiver5_irq                                          : std_logic;                      -- dma_dconvi:dma_ctl_irq -> irq_mapper_001:receiver5_irq
	signal irq_mapper_001_receiver6_irq                                          : std_logic;                      -- dma_dconvq:dma_ctl_irq -> irq_mapper_001:receiver6_irq
	signal irq_mapper_001_receiver7_irq                                          : std_logic;                      -- spi_afe_relays:irq -> irq_mapper_001:receiver7_irq
	signal hps_0_f2h_irq1_irq                                                    : std_logic_vector(31 downto 0);  -- irq_mapper_001:sender_irq -> hps_0:f2h_irq_p1
	signal adc_fifo_dc_out_valid                                                 : std_logic;                      -- adc_fifo_dc:out_valid -> avalon_st_adapter:in_0_valid
	signal adc_fifo_dc_out_data                                                  : std_logic_vector(15 downto 0);  -- adc_fifo_dc:out_data -> avalon_st_adapter:in_0_data
	signal adc_fifo_dc_out_ready                                                 : std_logic;                      -- avalon_st_adapter:in_0_ready -> adc_fifo_dc:out_ready
	signal avalon_st_adapter_out_0_valid                                         : std_logic;                      -- avalon_st_adapter:out_0_valid -> adc_fifo_mem:avalonst_sink_valid
	signal avalon_st_adapter_out_0_data                                          : std_logic_vector(31 downto 0);  -- avalon_st_adapter:out_0_data -> adc_fifo_mem:avalonst_sink_data
	signal avalon_st_adapter_out_0_ready                                         : std_logic;                      -- adc_fifo_mem:avalonst_sink_ready -> avalon_st_adapter:out_0_ready
	signal dconv_fifo_dc_out_valid                                               : std_logic;                      -- dconv_fifo_dc:out_valid -> avalon_st_adapter_001:in_0_valid
	signal dconv_fifo_dc_out_data                                                : std_logic_vector(31 downto 0);  -- dconv_fifo_dc:out_data -> avalon_st_adapter_001:in_0_data
	signal dconv_fifo_dc_out_ready                                               : std_logic;                      -- avalon_st_adapter_001:in_0_ready -> dconv_fifo_dc:out_ready
	signal avalon_st_adapter_001_out_0_valid                                     : std_logic;                      -- avalon_st_adapter_001:out_0_valid -> dconv_fifo_mem:avalonst_sink_valid
	signal avalon_st_adapter_001_out_0_data                                      : std_logic_vector(31 downto 0);  -- avalon_st_adapter_001:out_0_data -> dconv_fifo_mem:avalonst_sink_data
	signal avalon_st_adapter_001_out_0_ready                                     : std_logic;                      -- dconv_fifo_mem:avalonst_sink_ready -> avalon_st_adapter_001:out_0_ready
	signal dconv_fifo_dc_q_out_valid                                             : std_logic;                      -- dconv_fifo_dc_q:out_valid -> avalon_st_adapter_002:in_0_valid
	signal dconv_fifo_dc_q_out_data                                              : std_logic_vector(31 downto 0);  -- dconv_fifo_dc_q:out_data -> avalon_st_adapter_002:in_0_data
	signal dconv_fifo_dc_q_out_ready                                             : std_logic;                      -- avalon_st_adapter_002:in_0_ready -> dconv_fifo_dc_q:out_ready
	signal avalon_st_adapter_002_out_0_valid                                     : std_logic;                      -- avalon_st_adapter_002:out_0_valid -> dconv_fifo_mem_q:avalonst_sink_valid
	signal avalon_st_adapter_002_out_0_data                                      : std_logic_vector(31 downto 0);  -- avalon_st_adapter_002:out_0_data -> dconv_fifo_mem_q:avalonst_sink_data
	signal avalon_st_adapter_002_out_0_ready                                     : std_logic;                      -- dconv_fifo_mem_q:avalonst_sink_ready -> avalon_st_adapter_002:out_0_ready
	signal rst_controller_reset_out_reset                                        : std_logic;                      -- rst_controller:reset_out -> rst_controller_reset_out_reset:in
	signal rst_controller_001_reset_out_reset                                    : std_logic;                      -- rst_controller_001:reset_out -> [avalon_st_adapter:in_rst_0_reset, avalon_st_adapter_001:in_rst_0_reset, avalon_st_adapter_002:in_rst_0_reset, mm_interconnect_1:adc_fifo_mem_reset_in_reset_bridge_in_reset_reset, rst_controller_001_reset_out_reset:in]
	signal rst_controller_002_reset_out_reset                                    : std_logic;                      -- rst_controller_002:reset_out -> [alt_vip_itc_0:rst, alt_vip_vfr_vga:reset, mm_interconnect_1:alt_vip_vfr_vga_clock_reset_reset_reset_bridge_in_reset_reset]
	signal rst_controller_003_reset_out_reset                                    : std_logic;                      -- rst_controller_003:reset_out -> [alt_vip_vfr_vga:master_reset, analyzer_pll_reconfig:mgmt_reset, mm_interconnect_0:alt_vip_vfr_vga_clock_master_reset_reset_bridge_in_reset_reset, mm_interconnect_0:master_secure_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_1:dma_fifo_reset_reset_bridge_in_reset_reset, mm_interconnect_1:master_non_sec_clk_reset_reset_bridge_in_reset_reset, nmr_sys_pll_reconfig:mgmt_reset, rst_controller_003_reset_out_reset:in]
	signal rst_controller_004_reset_out_reset                                    : std_logic;                      -- rst_controller_004:reset_out -> [mm_interconnect_0:hps_0_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_1:hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset]
	signal fifo_rst_reset_ports_inv                                              : std_logic;                      -- fifo_rst_reset:inv -> [dconv_fir:reset_n, dconv_fir_q:reset_n]
	signal hps_0_h2f_reset_reset_n_ports_inv                                     : std_logic;                      -- hps_0_h2f_reset_reset_n:inv -> rst_controller_004:reset_in0
	signal reset_reset_n_ports_inv                                               : std_logic;                      -- reset_reset_n:inv -> [gp_pll:rst, master_non_sec:clk_reset_reset, master_secure:clk_reset_reset, rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_002:reset_in0, rst_controller_003:reset_in0]
	signal dma_fifo_write_master_write_ports_inv                                 : std_logic;                      -- dma_fifo_write_master_write:inv -> mm_interconnect_1:dma_fifo_write_master_write
	signal dma_dconvi_write_master_write_ports_inv                               : std_logic;                      -- dma_dconvi_write_master_write:inv -> mm_interconnect_1:dma_dconvi_write_master_write
	signal dma_dconvq_write_master_write_ports_inv                               : std_logic;                      -- dma_dconvq_write_master_write:inv -> mm_interconnect_1:dma_dconvq_write_master_write
	signal dma_dummy_write_master_write_ports_inv                                : std_logic;                      -- dma_dummy_write_master_write:inv -> mm_interconnect_1:dma_dummy_write_master_write
	signal dma_fifo_read_master_read_ports_inv                                   : std_logic;                      -- dma_fifo_read_master_read:inv -> mm_interconnect_1:dma_fifo_read_master_read
	signal dma_dconvq_read_master_read_ports_inv                                 : std_logic;                      -- dma_dconvq_read_master_read:inv -> mm_interconnect_1:dma_dconvq_read_master_read
	signal dma_dconvi_read_master_read_ports_inv                                 : std_logic;                      -- dma_dconvi_read_master_read:inv -> mm_interconnect_1:dma_dconvi_read_master_read
	signal dma_dummy_read_master_read_ports_inv                                  : std_logic;                      -- dma_dummy_read_master_read:inv -> mm_interconnect_1:dma_dummy_read_master_read
	signal mm_interconnect_1_sdram_s1_read_ports_inv                             : std_logic;                      -- mm_interconnect_1_sdram_s1_read:inv -> sdram:az_rd_n
	signal mm_interconnect_1_sdram_s1_byteenable_ports_inv                       : std_logic_vector(1 downto 0);   -- mm_interconnect_1_sdram_s1_byteenable:inv -> sdram:az_be_n
	signal mm_interconnect_1_sdram_s1_write_ports_inv                            : std_logic;                      -- mm_interconnect_1_sdram_s1_write:inv -> sdram:az_wr_n
	signal mm_interconnect_1_nmr_parameters_adc_val_sub_s1_write_ports_inv       : std_logic;                      -- mm_interconnect_1_nmr_parameters_adc_val_sub_s1_write:inv -> nmr_parameters:adc_val_sub_s1_write_n
	signal mm_interconnect_1_jtag_uart_avalon_jtag_slave_read_ports_inv          : std_logic;                      -- mm_interconnect_1_jtag_uart_avalon_jtag_slave_read:inv -> jtag_uart:av_read_n
	signal mm_interconnect_1_jtag_uart_avalon_jtag_slave_write_ports_inv         : std_logic;                      -- mm_interconnect_1_jtag_uart_avalon_jtag_slave_write:inv -> jtag_uart:av_write_n
	signal mm_interconnect_1_nmr_parameters_delay_nosig_s1_write_ports_inv       : std_logic;                      -- mm_interconnect_1_nmr_parameters_delay_nosig_s1_write:inv -> nmr_parameters:delay_nosig_s1_write_n
	signal mm_interconnect_1_nmr_parameters_delay_sig_s1_write_ports_inv         : std_logic;                      -- mm_interconnect_1_nmr_parameters_delay_sig_s1_write:inv -> nmr_parameters:delay_sig_s1_write_n
	signal mm_interconnect_1_nmr_parameters_delay_t1_s1_write_ports_inv          : std_logic;                      -- mm_interconnect_1_nmr_parameters_delay_t1_s1_write:inv -> nmr_parameters:delay_t1_s1_write_n
	signal mm_interconnect_1_nmr_parameters_echoes_per_scan_s1_write_ports_inv   : std_logic;                      -- mm_interconnect_1_nmr_parameters_echoes_per_scan_s1_write:inv -> nmr_parameters:echoes_per_scan_s1_write_n
	signal mm_interconnect_1_nmr_parameters_init_delay_s1_write_ports_inv        : std_logic;                      -- mm_interconnect_1_nmr_parameters_init_delay_s1_write:inv -> nmr_parameters:init_delay_s1_write_n
	signal mm_interconnect_1_nmr_parameters_pulse_180deg_s1_write_ports_inv      : std_logic;                      -- mm_interconnect_1_nmr_parameters_pulse_180deg_s1_write:inv -> nmr_parameters:pulse_180deg_s1_write_n
	signal mm_interconnect_1_nmr_parameters_pulse_90deg_s1_write_ports_inv       : std_logic;                      -- mm_interconnect_1_nmr_parameters_pulse_90deg_s1_write:inv -> nmr_parameters:pulse_90deg_s1_write_n
	signal mm_interconnect_1_nmr_parameters_pulse_t1_s1_write_ports_inv          : std_logic;                      -- mm_interconnect_1_nmr_parameters_pulse_t1_s1_write:inv -> nmr_parameters:pulse_t1_s1_write_n
	signal mm_interconnect_1_nmr_parameters_rx_delay_s1_write_ports_inv          : std_logic;                      -- mm_interconnect_1_nmr_parameters_rx_delay_s1_write:inv -> nmr_parameters:rx_delay_s1_write_n
	signal mm_interconnect_1_ctrl_out_s1_write_ports_inv                         : std_logic;                      -- mm_interconnect_1_ctrl_out_s1_write:inv -> ctrl_out:write_n
	signal mm_interconnect_1_aux_cnt_out_s1_write_ports_inv                      : std_logic;                      -- mm_interconnect_1_aux_cnt_out_s1_write:inv -> aux_cnt_out:write_n
	signal mm_interconnect_1_nmr_parameters_samples_per_echo_s1_write_ports_inv  : std_logic;                      -- mm_interconnect_1_nmr_parameters_samples_per_echo_s1_write:inv -> nmr_parameters:samples_per_echo_s1_write_n
	signal mm_interconnect_1_dac_grad_spi_control_port_read_ports_inv            : std_logic;                      -- mm_interconnect_1_dac_grad_spi_control_port_read:inv -> dac_grad:read_n
	signal mm_interconnect_1_dac_grad_spi_control_port_write_ports_inv           : std_logic;                      -- mm_interconnect_1_dac_grad_spi_control_port_write:inv -> dac_grad:write_n
	signal mm_interconnect_1_spi_mtch_ntwrk_spi_control_port_read_ports_inv      : std_logic;                      -- mm_interconnect_1_spi_mtch_ntwrk_spi_control_port_read:inv -> spi_mtch_ntwrk:read_n
	signal mm_interconnect_1_spi_mtch_ntwrk_spi_control_port_write_ports_inv     : std_logic;                      -- mm_interconnect_1_spi_mtch_ntwrk_spi_control_port_write:inv -> spi_mtch_ntwrk:write_n
	signal mm_interconnect_1_spi_afe_relays_spi_control_port_read_ports_inv      : std_logic;                      -- mm_interconnect_1_spi_afe_relays_spi_control_port_read:inv -> spi_afe_relays:read_n
	signal mm_interconnect_1_spi_afe_relays_spi_control_port_write_ports_inv     : std_logic;                      -- mm_interconnect_1_spi_afe_relays_spi_control_port_write:inv -> spi_afe_relays:write_n
	signal mm_interconnect_1_dma_fifo_control_port_slave_write_ports_inv         : std_logic;                      -- mm_interconnect_1_dma_fifo_control_port_slave_write:inv -> dma_fifo:dma_ctl_write_n
	signal mm_interconnect_1_dma_dconvi_control_port_slave_write_ports_inv       : std_logic;                      -- mm_interconnect_1_dma_dconvi_control_port_slave_write:inv -> dma_dconvi:dma_ctl_write_n
	signal mm_interconnect_1_dma_dconvq_control_port_slave_write_ports_inv       : std_logic;                      -- mm_interconnect_1_dma_dconvq_control_port_slave_write:inv -> dma_dconvq:dma_ctl_write_n
	signal mm_interconnect_1_dma_dummy_control_port_slave_write_ports_inv        : std_logic;                      -- mm_interconnect_1_dma_dummy_control_port_slave_write:inv -> dma_dummy:dma_ctl_write_n
	signal rst_controller_reset_out_reset_ports_inv                              : std_logic;                      -- rst_controller_reset_out_reset:inv -> [adc_fifo_dc:in_reset_n, dconv_fifo_dc:in_reset_n, dconv_fifo_dc_q:in_reset_n]
	signal rst_controller_001_reset_out_reset_ports_inv                          : std_logic;                      -- rst_controller_001_reset_out_reset:inv -> [adc_fifo_dc:out_reset_n, adc_fifo_mem:reset_n, dconv_fifo_dc:out_reset_n, dconv_fifo_dc_q:out_reset_n, dconv_fifo_mem:reset_n, dconv_fifo_mem_q:reset_n]
	signal rst_controller_003_reset_out_reset_ports_inv                          : std_logic;                      -- rst_controller_003_reset_out_reset:inv -> [aux_cnt_out:reset_n, ctrl_in:reset_n, ctrl_out:reset_n, dac_grad:reset_n, dconv_fir:coeff_in_areset, dconv_fir_q:coeff_in_areset, dma_dconvi:system_reset_n, dma_dconvq:system_reset_n, dma_dummy:system_reset_n, dma_fifo:system_reset_n, fifo_dummy64_in:reset_n, fifo_dummy64_out:reset_n, fifo_dummy:reset_n, i2c_ext:rst_n, i2c_int:rst_n, jtag_uart:rst_n, nmr_parameters:adc_val_sub_reset_reset_n, nmr_parameters:delay_nosig_reset_reset_n, nmr_parameters:delay_sig_reset_reset_n, nmr_parameters:delay_t1_reset_reset_n, nmr_parameters:echoes_per_scan_reset_reset_n, nmr_parameters:init_delay_reset_reset_n, nmr_parameters:pulse_180deg_reset_reset_n, nmr_parameters:pulse_90deg_reset_reset_n, nmr_parameters:pulse_t1_reset_reset_n, nmr_parameters:rx_delay_reset_reset_n, nmr_parameters:samples_per_echo_reset_reset_n, sdram:reset_n, spi_afe_relays:reset_n, spi_mtch_ntwrk:reset_n, switches:reset_n, sysid_qsys:reset_n]

begin

	adc_fifo_dc : component soc_system_v5_adc_fifo_dc
		generic map (
			SYMBOLS_PER_BEAT   => 1,
			BITS_PER_SYMBOL    => 16,
			FIFO_DEPTH         => 16384,
			CHANNEL_WIDTH      => 0,
			ERROR_WIDTH        => 0,
			USE_PACKETS        => 0,
			USE_IN_FILL_LEVEL  => 0,
			USE_OUT_FILL_LEVEL => 0,
			WR_SYNC_DEPTH      => 3,
			RD_SYNC_DEPTH      => 3
		)
		port map (
			in_clk            => fifo_clk_bridge_in_clk,                       --        in_clk.clk
			in_reset_n        => rst_controller_reset_out_reset_ports_inv,     --  in_clk_reset.reset_n
			out_clk           => clk_clk,                                      --       out_clk.clk
			out_reset_n       => rst_controller_001_reset_out_reset_ports_inv, -- out_clk_reset.reset_n
			in_data           => adc_fifo_in_data,                             --            in.data
			in_valid          => adc_fifo_in_valid,                            --              .valid
			in_ready          => adc_fifo_in_ready,                            --              .ready
			out_data          => adc_fifo_dc_out_data,                         --           out.data
			out_valid         => adc_fifo_dc_out_valid,                        --              .valid
			out_ready         => adc_fifo_dc_out_ready,                        --              .ready
			in_csr_address    => '0',                                          --   (terminated)
			in_csr_read       => '0',                                          --   (terminated)
			in_csr_write      => '0',                                          --   (terminated)
			in_csr_readdata   => open,                                         --   (terminated)
			in_csr_writedata  => "00000000000000000000000000000000",           --   (terminated)
			out_csr_address   => '0',                                          --   (terminated)
			out_csr_read      => '0',                                          --   (terminated)
			out_csr_write     => '0',                                          --   (terminated)
			out_csr_readdata  => open,                                         --   (terminated)
			out_csr_writedata => "00000000000000000000000000000000",           --   (terminated)
			in_startofpacket  => '0',                                          --   (terminated)
			in_endofpacket    => '0',                                          --   (terminated)
			out_startofpacket => open,                                         --   (terminated)
			out_endofpacket   => open,                                         --   (terminated)
			in_empty          => "0",                                          --   (terminated)
			out_empty         => open,                                         --   (terminated)
			in_error          => "0",                                          --   (terminated)
			out_error         => open,                                         --   (terminated)
			in_channel        => "0",                                          --   (terminated)
			out_channel       => open,                                         --   (terminated)
			space_avail_data  => open                                          --   (terminated)
		);

	adc_fifo_mem : component soc_system_v5_adc_fifo_mem
		port map (
			wrclock                         => clk_clk,                                         --   clk_in.clk
			reset_n                         => rst_controller_001_reset_out_reset_ports_inv,    -- reset_in.reset_n
			avalonst_sink_valid             => avalon_st_adapter_out_0_valid,                   --       in.valid
			avalonst_sink_data              => avalon_st_adapter_out_0_data,                    --         .data
			avalonst_sink_ready             => avalon_st_adapter_out_0_ready,                   --         .ready
			avalonmm_read_slave_readdata    => mm_interconnect_1_adc_fifo_mem_out_readdata,     --      out.readdata
			avalonmm_read_slave_read        => mm_interconnect_1_adc_fifo_mem_out_read,         --         .read
			avalonmm_read_slave_address     => mm_interconnect_1_adc_fifo_mem_out_address(0),   --         .address
			avalonmm_read_slave_waitrequest => mm_interconnect_1_adc_fifo_mem_out_waitrequest,  --         .waitrequest
			wrclk_control_slave_address     => mm_interconnect_1_adc_fifo_mem_in_csr_address,   --   in_csr.address
			wrclk_control_slave_read        => mm_interconnect_1_adc_fifo_mem_in_csr_read,      --         .read
			wrclk_control_slave_writedata   => mm_interconnect_1_adc_fifo_mem_in_csr_writedata, --         .writedata
			wrclk_control_slave_write       => mm_interconnect_1_adc_fifo_mem_in_csr_write,     --         .write
			wrclk_control_slave_readdata    => mm_interconnect_1_adc_fifo_mem_in_csr_readdata   --         .readdata
		);

	alt_vip_itc_0 : component soc_system_v5_alt_vip_itc_0
		port map (
			is_clk        => gp_pll_outclk0_clk,                                    --       is_clk_rst.clk
			rst           => rst_controller_002_reset_out_reset,                    -- is_clk_rst_reset.reset
			is_data       => alt_vip_vfr_vga_avalon_streaming_source_data,          --              din.data
			is_valid      => alt_vip_vfr_vga_avalon_streaming_source_valid,         --                 .valid
			is_ready      => alt_vip_vfr_vga_avalon_streaming_source_ready,         --                 .ready
			is_sop        => alt_vip_vfr_vga_avalon_streaming_source_startofpacket, --                 .startofpacket
			is_eop        => alt_vip_vfr_vga_avalon_streaming_source_endofpacket,   --                 .endofpacket
			vid_clk       => alt_vip_itc_0_clocked_video_vid_clk,                   --    clocked_video.export
			vid_data      => alt_vip_itc_0_clocked_video_vid_data,                  --                 .export
			underflow     => alt_vip_itc_0_clocked_video_underflow,                 --                 .export
			vid_datavalid => alt_vip_itc_0_clocked_video_vid_datavalid,             --                 .export
			vid_v_sync    => alt_vip_itc_0_clocked_video_vid_v_sync,                --                 .export
			vid_h_sync    => alt_vip_itc_0_clocked_video_vid_h_sync,                --                 .export
			vid_f         => alt_vip_itc_0_clocked_video_vid_f,                     --                 .export
			vid_h         => alt_vip_itc_0_clocked_video_vid_h,                     --                 .export
			vid_v         => alt_vip_itc_0_clocked_video_vid_v                      --                 .export
		);

	alt_vip_vfr_vga : component soc_system_v5_alt_vip_vfr_vga
		port map (
			clock                => gp_pll_outclk0_clk,                                       --             clock_reset.clk
			reset                => rst_controller_002_reset_out_reset,                       --       clock_reset_reset.reset
			master_clock         => clk_clk,                                                  --            clock_master.clk
			master_reset         => rst_controller_003_reset_out_reset,                       --      clock_master_reset.reset
			slave_address        => mm_interconnect_1_alt_vip_vfr_vga_avalon_slave_address,   --            avalon_slave.address
			slave_write          => mm_interconnect_1_alt_vip_vfr_vga_avalon_slave_write,     --                        .write
			slave_writedata      => mm_interconnect_1_alt_vip_vfr_vga_avalon_slave_writedata, --                        .writedata
			slave_read           => mm_interconnect_1_alt_vip_vfr_vga_avalon_slave_read,      --                        .read
			slave_readdata       => mm_interconnect_1_alt_vip_vfr_vga_avalon_slave_readdata,  --                        .readdata
			slave_irq            => irq_mapper_receiver0_irq,                                 --        interrupt_sender.irq
			dout_data            => alt_vip_vfr_vga_avalon_streaming_source_data,             -- avalon_streaming_source.data
			dout_valid           => alt_vip_vfr_vga_avalon_streaming_source_valid,            --                        .valid
			dout_ready           => alt_vip_vfr_vga_avalon_streaming_source_ready,            --                        .ready
			dout_startofpacket   => alt_vip_vfr_vga_avalon_streaming_source_startofpacket,    --                        .startofpacket
			dout_endofpacket     => alt_vip_vfr_vga_avalon_streaming_source_endofpacket,      --                        .endofpacket
			master_address       => alt_vip_vfr_vga_avalon_master_address,                    --           avalon_master.address
			master_burstcount    => alt_vip_vfr_vga_avalon_master_burstcount,                 --                        .burstcount
			master_readdata      => alt_vip_vfr_vga_avalon_master_readdata,                   --                        .readdata
			master_read          => alt_vip_vfr_vga_avalon_master_read,                       --                        .read
			master_readdatavalid => alt_vip_vfr_vga_avalon_master_readdatavalid,              --                        .readdatavalid
			master_waitrequest   => alt_vip_vfr_vga_avalon_master_waitrequest                 --                        .waitrequest
		);

	analyzer_pll : component soc_system_v5_analyzer_pll
		port map (
			refclk            => clk_clk,                                               --            refclk.clk
			rst               => analyzer_pll_reset_reset,                              --             reset.reset
			outclk_0          => analyzer_pll_outclk0_clk,                              --           outclk0.clk
			outclk_1          => analyzer_pll_outclk1_clk,                              --           outclk1.clk
			outclk_2          => analyzer_pll_outclk2_clk,                              --           outclk2.clk
			outclk_3          => analyzer_pll_outclk3_clk,                              --           outclk3.clk
			locked            => analyzer_pll_locked_export,                            --            locked.export
			reconfig_to_pll   => analyzer_pll_reconfig_reconfig_to_pll_reconfig_to_pll, --   reconfig_to_pll.reconfig_to_pll
			reconfig_from_pll => analyzer_pll_reconfig_from_pll_reconfig_from_pll       -- reconfig_from_pll.reconfig_from_pll
		);

	analyzer_pll_reconfig : component altera_pll_reconfig_top
		generic map (
			device_family       => "Cyclone V",
			ENABLE_MIF          => false,
			MIF_FILE_NAME       => "",
			ENABLE_BYTEENABLE   => false,
			BYTEENABLE_WIDTH    => 4,
			RECONFIG_ADDR_WIDTH => 6,
			RECONFIG_DATA_WIDTH => 32,
			reconf_width        => 64,
			WAIT_FOR_LOCK       => true
		)
		port map (
			mgmt_clk          => clk_clk,                                                               --          mgmt_clk.clk
			mgmt_reset        => rst_controller_003_reset_out_reset,                                    --        mgmt_reset.reset
			mgmt_waitrequest  => mm_interconnect_1_analyzer_pll_reconfig_mgmt_avalon_slave_waitrequest, -- mgmt_avalon_slave.waitrequest
			mgmt_read         => mm_interconnect_1_analyzer_pll_reconfig_mgmt_avalon_slave_read,        --                  .read
			mgmt_write        => mm_interconnect_1_analyzer_pll_reconfig_mgmt_avalon_slave_write,       --                  .write
			mgmt_readdata     => mm_interconnect_1_analyzer_pll_reconfig_mgmt_avalon_slave_readdata,    --                  .readdata
			mgmt_address      => mm_interconnect_1_analyzer_pll_reconfig_mgmt_avalon_slave_address,     --                  .address
			mgmt_writedata    => mm_interconnect_1_analyzer_pll_reconfig_mgmt_avalon_slave_writedata,   --                  .writedata
			reconfig_to_pll   => analyzer_pll_reconfig_reconfig_to_pll_reconfig_to_pll,                 --   reconfig_to_pll.reconfig_to_pll
			reconfig_from_pll => analyzer_pll_reconfig_from_pll_reconfig_from_pll,                      -- reconfig_from_pll.reconfig_from_pll
			mgmt_byteenable   => "0000"                                                                 --       (terminated)
		);

	aux_cnt_out : component soc_system_v5_aux_cnt_out
		port map (
			clk        => clk_clk,                                          --                 clk.clk
			reset_n    => rst_controller_003_reset_out_reset_ports_inv,     --               reset.reset_n
			address    => mm_interconnect_1_aux_cnt_out_s1_address,         --                  s1.address
			write_n    => mm_interconnect_1_aux_cnt_out_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_1_aux_cnt_out_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_1_aux_cnt_out_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_1_aux_cnt_out_s1_readdata,        --                    .readdata
			out_port   => aux_cnt_out_export                                -- external_connection.export
		);

	ctrl_in : component soc_system_v5_ctrl_in
		port map (
			clk      => clk_clk,                                      --                 clk.clk
			reset_n  => rst_controller_003_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_1_ctrl_in_s1_address,         --                  s1.address
			readdata => mm_interconnect_1_ctrl_in_s1_readdata,        --                    .readdata
			in_port  => ctrl_in_export                                -- external_connection.export
		);

	ctrl_out : component soc_system_v5_aux_cnt_out
		port map (
			clk        => clk_clk,                                       --                 clk.clk
			reset_n    => rst_controller_003_reset_out_reset_ports_inv,  --               reset.reset_n
			address    => mm_interconnect_1_ctrl_out_s1_address,         --                  s1.address
			write_n    => mm_interconnect_1_ctrl_out_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_1_ctrl_out_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_1_ctrl_out_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_1_ctrl_out_s1_readdata,        --                    .readdata
			out_port   => ctrl_out_export                                -- external_connection.export
		);

	dac_grad : component soc_system_v5_dac_grad
		port map (
			clk           => clk_clk,                                                     --              clk.clk
			reset_n       => rst_controller_003_reset_out_reset_ports_inv,                --            reset.reset_n
			data_from_cpu => mm_interconnect_1_dac_grad_spi_control_port_writedata,       -- spi_control_port.writedata
			data_to_cpu   => mm_interconnect_1_dac_grad_spi_control_port_readdata,        --                 .readdata
			mem_addr      => mm_interconnect_1_dac_grad_spi_control_port_address,         --                 .address
			read_n        => mm_interconnect_1_dac_grad_spi_control_port_read_ports_inv,  --                 .read_n
			spi_select    => mm_interconnect_1_dac_grad_spi_control_port_chipselect,      --                 .chipselect
			write_n       => mm_interconnect_1_dac_grad_spi_control_port_write_ports_inv, --                 .write_n
			irq           => irq_mapper_001_receiver2_irq,                                --              irq.irq
			MISO          => dac_grad_MISO,                                               --         external.export
			MOSI          => dac_grad_MOSI,                                               --                 .export
			SCLK          => dac_grad_SCLK,                                               --                 .export
			SS_n          => dac_grad_SS_n                                                --                 .export
		);

	dconv_fifo_dc : component soc_system_v5_dconv_fifo_dc
		generic map (
			SYMBOLS_PER_BEAT   => 1,
			BITS_PER_SYMBOL    => 32,
			FIFO_DEPTH         => 32768,
			CHANNEL_WIDTH      => 0,
			ERROR_WIDTH        => 0,
			USE_PACKETS        => 0,
			USE_IN_FILL_LEVEL  => 0,
			USE_OUT_FILL_LEVEL => 0,
			WR_SYNC_DEPTH      => 3,
			RD_SYNC_DEPTH      => 3
		)
		port map (
			in_clk            => fifo_clk_bridge_in_clk,                       --        in_clk.clk
			in_reset_n        => rst_controller_reset_out_reset_ports_inv,     --  in_clk_reset.reset_n
			out_clk           => clk_clk,                                      --       out_clk.clk
			out_reset_n       => rst_controller_001_reset_out_reset_ports_inv, -- out_clk_reset.reset_n
			in_data           => dconv_fifo_in_data,                           --            in.data
			in_valid          => dconv_fifo_in_valid,                          --              .valid
			in_ready          => dconv_fifo_in_ready,                          --              .ready
			out_data          => dconv_fifo_dc_out_data,                       --           out.data
			out_valid         => dconv_fifo_dc_out_valid,                      --              .valid
			out_ready         => dconv_fifo_dc_out_ready,                      --              .ready
			in_csr_address    => '0',                                          --   (terminated)
			in_csr_read       => '0',                                          --   (terminated)
			in_csr_write      => '0',                                          --   (terminated)
			in_csr_readdata   => open,                                         --   (terminated)
			in_csr_writedata  => "00000000000000000000000000000000",           --   (terminated)
			out_csr_address   => '0',                                          --   (terminated)
			out_csr_read      => '0',                                          --   (terminated)
			out_csr_write     => '0',                                          --   (terminated)
			out_csr_readdata  => open,                                         --   (terminated)
			out_csr_writedata => "00000000000000000000000000000000",           --   (terminated)
			in_startofpacket  => '0',                                          --   (terminated)
			in_endofpacket    => '0',                                          --   (terminated)
			out_startofpacket => open,                                         --   (terminated)
			out_endofpacket   => open,                                         --   (terminated)
			in_empty          => "0",                                          --   (terminated)
			out_empty         => open,                                         --   (terminated)
			in_error          => "0",                                          --   (terminated)
			out_error         => open,                                         --   (terminated)
			in_channel        => "0",                                          --   (terminated)
			out_channel       => open,                                         --   (terminated)
			space_avail_data  => open                                          --   (terminated)
		);

	dconv_fifo_dc_q : component soc_system_v5_dconv_fifo_dc
		generic map (
			SYMBOLS_PER_BEAT   => 1,
			BITS_PER_SYMBOL    => 32,
			FIFO_DEPTH         => 32768,
			CHANNEL_WIDTH      => 0,
			ERROR_WIDTH        => 0,
			USE_PACKETS        => 0,
			USE_IN_FILL_LEVEL  => 0,
			USE_OUT_FILL_LEVEL => 0,
			WR_SYNC_DEPTH      => 3,
			RD_SYNC_DEPTH      => 3
		)
		port map (
			in_clk            => fifo_clk_bridge_in_clk,                       --        in_clk.clk
			in_reset_n        => rst_controller_reset_out_reset_ports_inv,     --  in_clk_reset.reset_n
			out_clk           => clk_clk,                                      --       out_clk.clk
			out_reset_n       => rst_controller_001_reset_out_reset_ports_inv, -- out_clk_reset.reset_n
			in_data           => dconv_fifo_q_in_data,                         --            in.data
			in_valid          => dconv_fifo_q_in_valid,                        --              .valid
			in_ready          => dconv_fifo_q_in_ready,                        --              .ready
			out_data          => dconv_fifo_dc_q_out_data,                     --           out.data
			out_valid         => dconv_fifo_dc_q_out_valid,                    --              .valid
			out_ready         => dconv_fifo_dc_q_out_ready,                    --              .ready
			in_csr_address    => '0',                                          --   (terminated)
			in_csr_read       => '0',                                          --   (terminated)
			in_csr_write      => '0',                                          --   (terminated)
			in_csr_readdata   => open,                                         --   (terminated)
			in_csr_writedata  => "00000000000000000000000000000000",           --   (terminated)
			out_csr_address   => '0',                                          --   (terminated)
			out_csr_read      => '0',                                          --   (terminated)
			out_csr_write     => '0',                                          --   (terminated)
			out_csr_readdata  => open,                                         --   (terminated)
			out_csr_writedata => "00000000000000000000000000000000",           --   (terminated)
			in_startofpacket  => '0',                                          --   (terminated)
			in_endofpacket    => '0',                                          --   (terminated)
			out_startofpacket => open,                                         --   (terminated)
			out_endofpacket   => open,                                         --   (terminated)
			in_empty          => "0",                                          --   (terminated)
			out_empty         => open,                                         --   (terminated)
			in_error          => "0",                                          --   (terminated)
			out_error         => open,                                         --   (terminated)
			in_channel        => "0",                                          --   (terminated)
			out_channel       => open,                                         --   (terminated)
			space_avail_data  => open                                          --   (terminated)
		);

	dconv_fifo_mem : component soc_system_v5_dconv_fifo_mem
		port map (
			wrclock                         => clk_clk,                                           --   clk_in.clk
			reset_n                         => rst_controller_001_reset_out_reset_ports_inv,      -- reset_in.reset_n
			avalonst_sink_valid             => avalon_st_adapter_001_out_0_valid,                 --       in.valid
			avalonst_sink_data              => avalon_st_adapter_001_out_0_data,                  --         .data
			avalonst_sink_ready             => avalon_st_adapter_001_out_0_ready,                 --         .ready
			avalonmm_read_slave_readdata    => mm_interconnect_1_dconv_fifo_mem_out_readdata,     --      out.readdata
			avalonmm_read_slave_read        => mm_interconnect_1_dconv_fifo_mem_out_read,         --         .read
			avalonmm_read_slave_address     => mm_interconnect_1_dconv_fifo_mem_out_address(0),   --         .address
			avalonmm_read_slave_waitrequest => mm_interconnect_1_dconv_fifo_mem_out_waitrequest,  --         .waitrequest
			wrclk_control_slave_address     => mm_interconnect_1_dconv_fifo_mem_in_csr_address,   --   in_csr.address
			wrclk_control_slave_read        => mm_interconnect_1_dconv_fifo_mem_in_csr_read,      --         .read
			wrclk_control_slave_writedata   => mm_interconnect_1_dconv_fifo_mem_in_csr_writedata, --         .writedata
			wrclk_control_slave_write       => mm_interconnect_1_dconv_fifo_mem_in_csr_write,     --         .write
			wrclk_control_slave_readdata    => mm_interconnect_1_dconv_fifo_mem_in_csr_readdata   --         .readdata
		);

	dconv_fifo_mem_q : component soc_system_v5_dconv_fifo_mem
		port map (
			wrclock                         => clk_clk,                                             --   clk_in.clk
			reset_n                         => rst_controller_001_reset_out_reset_ports_inv,        -- reset_in.reset_n
			avalonst_sink_valid             => avalon_st_adapter_002_out_0_valid,                   --       in.valid
			avalonst_sink_data              => avalon_st_adapter_002_out_0_data,                    --         .data
			avalonst_sink_ready             => avalon_st_adapter_002_out_0_ready,                   --         .ready
			avalonmm_read_slave_readdata    => mm_interconnect_1_dconv_fifo_mem_q_out_readdata,     --      out.readdata
			avalonmm_read_slave_read        => mm_interconnect_1_dconv_fifo_mem_q_out_read,         --         .read
			avalonmm_read_slave_address     => mm_interconnect_1_dconv_fifo_mem_q_out_address(0),   --         .address
			avalonmm_read_slave_waitrequest => mm_interconnect_1_dconv_fifo_mem_q_out_waitrequest,  --         .waitrequest
			wrclk_control_slave_address     => mm_interconnect_1_dconv_fifo_mem_q_in_csr_address,   --   in_csr.address
			wrclk_control_slave_read        => mm_interconnect_1_dconv_fifo_mem_q_in_csr_read,      --         .read
			wrclk_control_slave_writedata   => mm_interconnect_1_dconv_fifo_mem_q_in_csr_writedata, --         .writedata
			wrclk_control_slave_write       => mm_interconnect_1_dconv_fifo_mem_q_in_csr_write,     --         .write
			wrclk_control_slave_readdata    => mm_interconnect_1_dconv_fifo_mem_q_in_csr_readdata   --         .readdata
		);

	dconv_fir : component soc_system_v5_dconv_fir
		port map (
			clk                => fifo_clk_bridge_in_clk,                                    --                     clk.clk
			reset_n            => fifo_rst_reset_ports_inv,                                  --                     rst.reset_n
			ast_sink_data      => dconv_fir_in_data,                                         --   avalon_streaming_sink.data
			ast_sink_valid     => dconv_fir_in_valid,                                        --                        .valid
			ast_sink_error     => dconv_fir_in_error,                                        --                        .error
			ast_source_data    => dconv_fir_out_data,                                        -- avalon_streaming_source.data
			ast_source_valid   => dconv_fir_out_valid,                                       --                        .valid
			ast_source_error   => dconv_fir_out_error,                                       --                        .error
			coeff_in_clk       => clk_clk,                                                   --             coeff_clock.clk
			coeff_in_areset    => rst_controller_003_reset_out_reset_ports_inv,              --             coeff_reset.reset_n
			coeff_in_address   => mm_interconnect_1_dconv_fir_avalon_mm_slave_address,       --         avalon_mm_slave.address
			coeff_in_read      => mm_interconnect_1_dconv_fir_avalon_mm_slave_read,          --                        .read
			coeff_out_valid(0) => mm_interconnect_1_dconv_fir_avalon_mm_slave_readdatavalid, --                        .readdatavalid
			coeff_out_data     => mm_interconnect_1_dconv_fir_avalon_mm_slave_readdata,      --                        .readdata
			coeff_in_we(0)     => mm_interconnect_1_dconv_fir_avalon_mm_slave_write,         --                        .write
			coeff_in_data      => mm_interconnect_1_dconv_fir_avalon_mm_slave_writedata      --                        .writedata
		);

	dconv_fir_q : component soc_system_v5_dconv_fir
		port map (
			clk                => fifo_clk_bridge_in_clk,                                      --                     clk.clk
			reset_n            => fifo_rst_reset_ports_inv,                                    --                     rst.reset_n
			ast_sink_data      => dconv_fir_q_in_data,                                         --   avalon_streaming_sink.data
			ast_sink_valid     => dconv_fir_q_in_valid,                                        --                        .valid
			ast_sink_error     => dconv_fir_q_in_error,                                        --                        .error
			ast_source_data    => dconv_fir_q_out_data,                                        -- avalon_streaming_source.data
			ast_source_valid   => dconv_fir_q_out_valid,                                       --                        .valid
			ast_source_error   => dconv_fir_q_out_error,                                       --                        .error
			coeff_in_clk       => clk_clk,                                                     --             coeff_clock.clk
			coeff_in_areset    => rst_controller_003_reset_out_reset_ports_inv,                --             coeff_reset.reset_n
			coeff_in_address   => mm_interconnect_1_dconv_fir_q_avalon_mm_slave_address,       --         avalon_mm_slave.address
			coeff_in_read      => mm_interconnect_1_dconv_fir_q_avalon_mm_slave_read,          --                        .read
			coeff_out_valid(0) => mm_interconnect_1_dconv_fir_q_avalon_mm_slave_readdatavalid, --                        .readdatavalid
			coeff_out_data     => mm_interconnect_1_dconv_fir_q_avalon_mm_slave_readdata,      --                        .readdata
			coeff_in_we(0)     => mm_interconnect_1_dconv_fir_q_avalon_mm_slave_write,         --                        .write
			coeff_in_data      => mm_interconnect_1_dconv_fir_q_avalon_mm_slave_writedata      --                        .writedata
		);

	dma_dconvi : component soc_system_v5_dma_dconvi
		port map (
			clk                => clk_clk,                                                         --                clk.clk
			system_reset_n     => rst_controller_003_reset_out_reset_ports_inv,                    --              reset.reset_n
			dma_ctl_address    => mm_interconnect_1_dma_dconvi_control_port_slave_address,         -- control_port_slave.address
			dma_ctl_chipselect => mm_interconnect_1_dma_dconvi_control_port_slave_chipselect,      --                   .chipselect
			dma_ctl_readdata   => mm_interconnect_1_dma_dconvi_control_port_slave_readdata,        --                   .readdata
			dma_ctl_write_n    => mm_interconnect_1_dma_dconvi_control_port_slave_write_ports_inv, --                   .write_n
			dma_ctl_writedata  => mm_interconnect_1_dma_dconvi_control_port_slave_writedata,       --                   .writedata
			dma_ctl_irq        => irq_mapper_001_receiver5_irq,                                    --                irq.irq
			read_address       => dma_dconvi_read_master_address,                                  --        read_master.address
			read_chipselect    => dma_dconvi_read_master_chipselect,                               --                   .chipselect
			read_read_n        => dma_dconvi_read_master_read,                                     --                   .read_n
			read_readdata      => dma_dconvi_read_master_readdata,                                 --                   .readdata
			read_readdatavalid => dma_dconvi_read_master_readdatavalid,                            --                   .readdatavalid
			read_waitrequest   => dma_dconvi_read_master_waitrequest,                              --                   .waitrequest
			write_address      => dma_dconvi_write_master_address,                                 --       write_master.address
			write_chipselect   => dma_dconvi_write_master_chipselect,                              --                   .chipselect
			write_waitrequest  => dma_dconvi_write_master_waitrequest,                             --                   .waitrequest
			write_write_n      => dma_dconvi_write_master_write,                                   --                   .write_n
			write_writedata    => dma_dconvi_write_master_writedata,                               --                   .writedata
			write_byteenable   => dma_dconvi_write_master_byteenable                               --                   .byteenable
		);

	dma_dconvq : component soc_system_v5_dma_dconvq
		port map (
			clk                => clk_clk,                                                         --                clk.clk
			system_reset_n     => rst_controller_003_reset_out_reset_ports_inv,                    --              reset.reset_n
			dma_ctl_address    => mm_interconnect_1_dma_dconvq_control_port_slave_address,         -- control_port_slave.address
			dma_ctl_chipselect => mm_interconnect_1_dma_dconvq_control_port_slave_chipselect,      --                   .chipselect
			dma_ctl_readdata   => mm_interconnect_1_dma_dconvq_control_port_slave_readdata,        --                   .readdata
			dma_ctl_write_n    => mm_interconnect_1_dma_dconvq_control_port_slave_write_ports_inv, --                   .write_n
			dma_ctl_writedata  => mm_interconnect_1_dma_dconvq_control_port_slave_writedata,       --                   .writedata
			dma_ctl_irq        => irq_mapper_001_receiver6_irq,                                    --                irq.irq
			read_address       => dma_dconvq_read_master_address,                                  --        read_master.address
			read_chipselect    => dma_dconvq_read_master_chipselect,                               --                   .chipselect
			read_read_n        => dma_dconvq_read_master_read,                                     --                   .read_n
			read_readdata      => dma_dconvq_read_master_readdata,                                 --                   .readdata
			read_readdatavalid => dma_dconvq_read_master_readdatavalid,                            --                   .readdatavalid
			read_waitrequest   => dma_dconvq_read_master_waitrequest,                              --                   .waitrequest
			write_address      => dma_dconvq_write_master_address,                                 --       write_master.address
			write_chipselect   => dma_dconvq_write_master_chipselect,                              --                   .chipselect
			write_waitrequest  => dma_dconvq_write_master_waitrequest,                             --                   .waitrequest
			write_write_n      => dma_dconvq_write_master_write,                                   --                   .write_n
			write_writedata    => dma_dconvq_write_master_writedata,                               --                   .writedata
			write_byteenable   => dma_dconvq_write_master_byteenable                               --                   .byteenable
		);

	dma_dummy : component soc_system_v5_dma_dummy
		port map (
			clk                => clk_clk,                                                        --                clk.clk
			system_reset_n     => rst_controller_003_reset_out_reset_ports_inv,                   --              reset.reset_n
			dma_ctl_address    => mm_interconnect_1_dma_dummy_control_port_slave_address,         -- control_port_slave.address
			dma_ctl_chipselect => mm_interconnect_1_dma_dummy_control_port_slave_chipselect,      --                   .chipselect
			dma_ctl_readdata   => mm_interconnect_1_dma_dummy_control_port_slave_readdata,        --                   .readdata
			dma_ctl_write_n    => mm_interconnect_1_dma_dummy_control_port_slave_write_ports_inv, --                   .write_n
			dma_ctl_writedata  => mm_interconnect_1_dma_dummy_control_port_slave_writedata,       --                   .writedata
			dma_ctl_irq        => open,                                                           --                irq.irq
			read_address       => dma_dummy_read_master_address,                                  --        read_master.address
			read_chipselect    => dma_dummy_read_master_chipselect,                               --                   .chipselect
			read_read_n        => dma_dummy_read_master_read,                                     --                   .read_n
			read_readdata      => dma_dummy_read_master_readdata,                                 --                   .readdata
			read_readdatavalid => dma_dummy_read_master_readdatavalid,                            --                   .readdatavalid
			read_waitrequest   => dma_dummy_read_master_waitrequest,                              --                   .waitrequest
			write_address      => dma_dummy_write_master_address,                                 --       write_master.address
			write_chipselect   => dma_dummy_write_master_chipselect,                              --                   .chipselect
			write_waitrequest  => dma_dummy_write_master_waitrequest,                             --                   .waitrequest
			write_write_n      => dma_dummy_write_master_write,                                   --                   .write_n
			write_writedata    => dma_dummy_write_master_writedata,                               --                   .writedata
			write_byteenable   => dma_dummy_write_master_byteenable                               --                   .byteenable
		);

	dma_fifo : component soc_system_v5_dma_fifo
		port map (
			clk                => clk_clk,                                                       --                clk.clk
			system_reset_n     => rst_controller_003_reset_out_reset_ports_inv,                  --              reset.reset_n
			dma_ctl_address    => mm_interconnect_1_dma_fifo_control_port_slave_address,         -- control_port_slave.address
			dma_ctl_chipselect => mm_interconnect_1_dma_fifo_control_port_slave_chipselect,      --                   .chipselect
			dma_ctl_readdata   => mm_interconnect_1_dma_fifo_control_port_slave_readdata,        --                   .readdata
			dma_ctl_write_n    => mm_interconnect_1_dma_fifo_control_port_slave_write_ports_inv, --                   .write_n
			dma_ctl_writedata  => mm_interconnect_1_dma_fifo_control_port_slave_writedata,       --                   .writedata
			dma_ctl_irq        => irq_mapper_001_receiver3_irq,                                  --                irq.irq
			read_address       => dma_fifo_read_master_address,                                  --        read_master.address
			read_chipselect    => dma_fifo_read_master_chipselect,                               --                   .chipselect
			read_read_n        => dma_fifo_read_master_read,                                     --                   .read_n
			read_readdata      => dma_fifo_read_master_readdata,                                 --                   .readdata
			read_readdatavalid => dma_fifo_read_master_readdatavalid,                            --                   .readdatavalid
			read_waitrequest   => dma_fifo_read_master_waitrequest,                              --                   .waitrequest
			write_address      => dma_fifo_write_master_address,                                 --       write_master.address
			write_chipselect   => dma_fifo_write_master_chipselect,                              --                   .chipselect
			write_waitrequest  => dma_fifo_write_master_waitrequest,                             --                   .waitrequest
			write_write_n      => dma_fifo_write_master_write,                                   --                   .write_n
			write_writedata    => dma_fifo_write_master_writedata,                               --                   .writedata
			write_byteenable   => dma_fifo_write_master_byteenable                               --                   .byteenable
		);

	fifo_dummy : component soc_system_v5_fifo_dummy
		port map (
			wrclock                          => clk_clk,                                       --   clk_in.clk
			reset_n                          => rst_controller_003_reset_out_reset_ports_inv,  -- reset_in.reset_n
			avalonmm_write_slave_writedata   => mm_interconnect_1_fifo_dummy_in_writedata,     --       in.writedata
			avalonmm_write_slave_write       => mm_interconnect_1_fifo_dummy_in_write,         --         .write
			avalonmm_write_slave_waitrequest => mm_interconnect_1_fifo_dummy_in_waitrequest,   --         .waitrequest
			avalonmm_read_slave_readdata     => mm_interconnect_1_fifo_dummy_out_readdata,     --      out.readdata
			avalonmm_read_slave_read         => mm_interconnect_1_fifo_dummy_out_read,         --         .read
			avalonmm_read_slave_waitrequest  => mm_interconnect_1_fifo_dummy_out_waitrequest,  --         .waitrequest
			wrclk_control_slave_address      => mm_interconnect_1_fifo_dummy_in_csr_address,   --   in_csr.address
			wrclk_control_slave_read         => mm_interconnect_1_fifo_dummy_in_csr_read,      --         .read
			wrclk_control_slave_writedata    => mm_interconnect_1_fifo_dummy_in_csr_writedata, --         .writedata
			wrclk_control_slave_write        => mm_interconnect_1_fifo_dummy_in_csr_write,     --         .write
			wrclk_control_slave_readdata     => mm_interconnect_1_fifo_dummy_in_csr_readdata   --         .readdata
		);

	fifo_dummy64_in : component soc_system_v5_fifo_dummy64_in
		port map (
			wrclock                          => clk_clk,                                            --   clk_in.clk
			reset_n                          => rst_controller_003_reset_out_reset_ports_inv,       -- reset_in.reset_n
			avalonmm_write_slave_writedata   => mm_interconnect_1_fifo_dummy64_in_in_writedata,     --       in.writedata
			avalonmm_write_slave_write       => mm_interconnect_1_fifo_dummy64_in_in_write,         --         .write
			avalonmm_write_slave_address     => mm_interconnect_1_fifo_dummy64_in_in_address(0),    --         .address
			avalonmm_write_slave_waitrequest => mm_interconnect_1_fifo_dummy64_in_in_waitrequest,   --         .waitrequest
			avalonst_source_valid            => fifo_dummy64_in_out_valid,                          --      out.valid
			avalonst_source_data             => fifo_dummy64_in_out_data,                           --         .data
			avalonst_source_ready            => fifo_dummy64_in_out_ready,                          --         .ready
			wrclk_control_slave_address      => mm_interconnect_1_fifo_dummy64_in_in_csr_address,   --   in_csr.address
			wrclk_control_slave_read         => mm_interconnect_1_fifo_dummy64_in_in_csr_read,      --         .read
			wrclk_control_slave_writedata    => mm_interconnect_1_fifo_dummy64_in_in_csr_writedata, --         .writedata
			wrclk_control_slave_write        => mm_interconnect_1_fifo_dummy64_in_in_csr_write,     --         .write
			wrclk_control_slave_readdata     => mm_interconnect_1_fifo_dummy64_in_in_csr_readdata   --         .readdata
		);

	fifo_dummy64_out : component soc_system_v5_fifo_dummy64_out
		port map (
			wrclock                         => clk_clk,                                             --   clk_in.clk
			reset_n                         => rst_controller_003_reset_out_reset_ports_inv,        -- reset_in.reset_n
			avalonst_sink_valid             => fifo_dummy64_in_out_valid,                           --       in.valid
			avalonst_sink_data              => fifo_dummy64_in_out_data,                            --         .data
			avalonst_sink_ready             => fifo_dummy64_in_out_ready,                           --         .ready
			avalonmm_read_slave_readdata    => mm_interconnect_1_fifo_dummy64_out_out_readdata,     --      out.readdata
			avalonmm_read_slave_read        => mm_interconnect_1_fifo_dummy64_out_out_read,         --         .read
			avalonmm_read_slave_address     => mm_interconnect_1_fifo_dummy64_out_out_address(0),   --         .address
			avalonmm_read_slave_waitrequest => mm_interconnect_1_fifo_dummy64_out_out_waitrequest,  --         .waitrequest
			wrclk_control_slave_address     => mm_interconnect_1_fifo_dummy64_out_in_csr_address,   --   in_csr.address
			wrclk_control_slave_read        => mm_interconnect_1_fifo_dummy64_out_in_csr_read,      --         .read
			wrclk_control_slave_writedata   => mm_interconnect_1_fifo_dummy64_out_in_csr_writedata, --         .writedata
			wrclk_control_slave_write       => mm_interconnect_1_fifo_dummy64_out_in_csr_write,     --         .write
			wrclk_control_slave_readdata    => mm_interconnect_1_fifo_dummy64_out_in_csr_readdata   --         .readdata
		);

	gp_pll : component soc_system_v5_gp_pll
		port map (
			refclk   => clk_clk,                 --  refclk.clk
			rst      => reset_reset_n_ports_inv, --   reset.reset
			outclk_0 => gp_pll_outclk0_clk,      -- outclk0.clk
			outclk_1 => pll_vga_clk65_clk,       -- outclk1.clk
			outclk_2 => open,                    -- outclk2.clk
			outclk_3 => sdram_clk_clk,           -- outclk3.clk
			locked   => pll_vga_locked_export    --  locked.export
		);

	hps_0 : component soc_system_v5_hps_0
		generic map (
			F2S_Width => 3,
			S2F_Width => 3
		)
		port map (
			mem_a                    => memory_mem_a,                                  --            memory.mem_a
			mem_ba                   => memory_mem_ba,                                 --                  .mem_ba
			mem_ck                   => memory_mem_ck,                                 --                  .mem_ck
			mem_ck_n                 => memory_mem_ck_n,                               --                  .mem_ck_n
			mem_cke                  => memory_mem_cke,                                --                  .mem_cke
			mem_cs_n                 => memory_mem_cs_n,                               --                  .mem_cs_n
			mem_ras_n                => memory_mem_ras_n,                              --                  .mem_ras_n
			mem_cas_n                => memory_mem_cas_n,                              --                  .mem_cas_n
			mem_we_n                 => memory_mem_we_n,                               --                  .mem_we_n
			mem_reset_n              => memory_mem_reset_n,                            --                  .mem_reset_n
			mem_dq                   => memory_mem_dq,                                 --                  .mem_dq
			mem_dqs                  => memory_mem_dqs,                                --                  .mem_dqs
			mem_dqs_n                => memory_mem_dqs_n,                              --                  .mem_dqs_n
			mem_odt                  => memory_mem_odt,                                --                  .mem_odt
			mem_dm                   => memory_mem_dm,                                 --                  .mem_dm
			oct_rzqin                => memory_oct_rzqin,                              --                  .oct_rzqin
			hps_io_emac1_inst_TX_CLK => hps_0_hps_io_hps_io_emac1_inst_TX_CLK,         --            hps_io.hps_io_emac1_inst_TX_CLK
			hps_io_emac1_inst_TXD0   => hps_0_hps_io_hps_io_emac1_inst_TXD0,           --                  .hps_io_emac1_inst_TXD0
			hps_io_emac1_inst_TXD1   => hps_0_hps_io_hps_io_emac1_inst_TXD1,           --                  .hps_io_emac1_inst_TXD1
			hps_io_emac1_inst_TXD2   => hps_0_hps_io_hps_io_emac1_inst_TXD2,           --                  .hps_io_emac1_inst_TXD2
			hps_io_emac1_inst_TXD3   => hps_0_hps_io_hps_io_emac1_inst_TXD3,           --                  .hps_io_emac1_inst_TXD3
			hps_io_emac1_inst_RXD0   => hps_0_hps_io_hps_io_emac1_inst_RXD0,           --                  .hps_io_emac1_inst_RXD0
			hps_io_emac1_inst_MDIO   => hps_0_hps_io_hps_io_emac1_inst_MDIO,           --                  .hps_io_emac1_inst_MDIO
			hps_io_emac1_inst_MDC    => hps_0_hps_io_hps_io_emac1_inst_MDC,            --                  .hps_io_emac1_inst_MDC
			hps_io_emac1_inst_RX_CTL => hps_0_hps_io_hps_io_emac1_inst_RX_CTL,         --                  .hps_io_emac1_inst_RX_CTL
			hps_io_emac1_inst_TX_CTL => hps_0_hps_io_hps_io_emac1_inst_TX_CTL,         --                  .hps_io_emac1_inst_TX_CTL
			hps_io_emac1_inst_RX_CLK => hps_0_hps_io_hps_io_emac1_inst_RX_CLK,         --                  .hps_io_emac1_inst_RX_CLK
			hps_io_emac1_inst_RXD1   => hps_0_hps_io_hps_io_emac1_inst_RXD1,           --                  .hps_io_emac1_inst_RXD1
			hps_io_emac1_inst_RXD2   => hps_0_hps_io_hps_io_emac1_inst_RXD2,           --                  .hps_io_emac1_inst_RXD2
			hps_io_emac1_inst_RXD3   => hps_0_hps_io_hps_io_emac1_inst_RXD3,           --                  .hps_io_emac1_inst_RXD3
			hps_io_qspi_inst_IO0     => hps_0_hps_io_hps_io_qspi_inst_IO0,             --                  .hps_io_qspi_inst_IO0
			hps_io_qspi_inst_IO1     => hps_0_hps_io_hps_io_qspi_inst_IO1,             --                  .hps_io_qspi_inst_IO1
			hps_io_qspi_inst_IO2     => hps_0_hps_io_hps_io_qspi_inst_IO2,             --                  .hps_io_qspi_inst_IO2
			hps_io_qspi_inst_IO3     => hps_0_hps_io_hps_io_qspi_inst_IO3,             --                  .hps_io_qspi_inst_IO3
			hps_io_qspi_inst_SS0     => hps_0_hps_io_hps_io_qspi_inst_SS0,             --                  .hps_io_qspi_inst_SS0
			hps_io_qspi_inst_CLK     => hps_0_hps_io_hps_io_qspi_inst_CLK,             --                  .hps_io_qspi_inst_CLK
			hps_io_sdio_inst_CMD     => hps_0_hps_io_hps_io_sdio_inst_CMD,             --                  .hps_io_sdio_inst_CMD
			hps_io_sdio_inst_D0      => hps_0_hps_io_hps_io_sdio_inst_D0,              --                  .hps_io_sdio_inst_D0
			hps_io_sdio_inst_D1      => hps_0_hps_io_hps_io_sdio_inst_D1,              --                  .hps_io_sdio_inst_D1
			hps_io_sdio_inst_CLK     => hps_0_hps_io_hps_io_sdio_inst_CLK,             --                  .hps_io_sdio_inst_CLK
			hps_io_sdio_inst_D2      => hps_0_hps_io_hps_io_sdio_inst_D2,              --                  .hps_io_sdio_inst_D2
			hps_io_sdio_inst_D3      => hps_0_hps_io_hps_io_sdio_inst_D3,              --                  .hps_io_sdio_inst_D3
			hps_io_usb1_inst_D0      => hps_0_hps_io_hps_io_usb1_inst_D0,              --                  .hps_io_usb1_inst_D0
			hps_io_usb1_inst_D1      => hps_0_hps_io_hps_io_usb1_inst_D1,              --                  .hps_io_usb1_inst_D1
			hps_io_usb1_inst_D2      => hps_0_hps_io_hps_io_usb1_inst_D2,              --                  .hps_io_usb1_inst_D2
			hps_io_usb1_inst_D3      => hps_0_hps_io_hps_io_usb1_inst_D3,              --                  .hps_io_usb1_inst_D3
			hps_io_usb1_inst_D4      => hps_0_hps_io_hps_io_usb1_inst_D4,              --                  .hps_io_usb1_inst_D4
			hps_io_usb1_inst_D5      => hps_0_hps_io_hps_io_usb1_inst_D5,              --                  .hps_io_usb1_inst_D5
			hps_io_usb1_inst_D6      => hps_0_hps_io_hps_io_usb1_inst_D6,              --                  .hps_io_usb1_inst_D6
			hps_io_usb1_inst_D7      => hps_0_hps_io_hps_io_usb1_inst_D7,              --                  .hps_io_usb1_inst_D7
			hps_io_usb1_inst_CLK     => hps_0_hps_io_hps_io_usb1_inst_CLK,             --                  .hps_io_usb1_inst_CLK
			hps_io_usb1_inst_STP     => hps_0_hps_io_hps_io_usb1_inst_STP,             --                  .hps_io_usb1_inst_STP
			hps_io_usb1_inst_DIR     => hps_0_hps_io_hps_io_usb1_inst_DIR,             --                  .hps_io_usb1_inst_DIR
			hps_io_usb1_inst_NXT     => hps_0_hps_io_hps_io_usb1_inst_NXT,             --                  .hps_io_usb1_inst_NXT
			hps_io_spim1_inst_CLK    => hps_0_hps_io_hps_io_spim1_inst_CLK,            --                  .hps_io_spim1_inst_CLK
			hps_io_spim1_inst_MOSI   => hps_0_hps_io_hps_io_spim1_inst_MOSI,           --                  .hps_io_spim1_inst_MOSI
			hps_io_spim1_inst_MISO   => hps_0_hps_io_hps_io_spim1_inst_MISO,           --                  .hps_io_spim1_inst_MISO
			hps_io_spim1_inst_SS0    => hps_0_hps_io_hps_io_spim1_inst_SS0,            --                  .hps_io_spim1_inst_SS0
			hps_io_uart0_inst_RX     => hps_0_hps_io_hps_io_uart0_inst_RX,             --                  .hps_io_uart0_inst_RX
			hps_io_uart0_inst_TX     => hps_0_hps_io_hps_io_uart0_inst_TX,             --                  .hps_io_uart0_inst_TX
			hps_io_i2c0_inst_SDA     => hps_0_hps_io_hps_io_i2c0_inst_SDA,             --                  .hps_io_i2c0_inst_SDA
			hps_io_i2c0_inst_SCL     => hps_0_hps_io_hps_io_i2c0_inst_SCL,             --                  .hps_io_i2c0_inst_SCL
			hps_io_i2c1_inst_SDA     => hps_0_hps_io_hps_io_i2c1_inst_SDA,             --                  .hps_io_i2c1_inst_SDA
			hps_io_i2c1_inst_SCL     => hps_0_hps_io_hps_io_i2c1_inst_SCL,             --                  .hps_io_i2c1_inst_SCL
			hps_io_gpio_inst_GPIO09  => hps_0_hps_io_hps_io_gpio_inst_GPIO09,          --                  .hps_io_gpio_inst_GPIO09
			hps_io_gpio_inst_GPIO35  => hps_0_hps_io_hps_io_gpio_inst_GPIO35,          --                  .hps_io_gpio_inst_GPIO35
			hps_io_gpio_inst_GPIO40  => hps_0_hps_io_hps_io_gpio_inst_GPIO40,          --                  .hps_io_gpio_inst_GPIO40
			hps_io_gpio_inst_GPIO48  => hps_0_hps_io_hps_io_gpio_inst_GPIO48,          --                  .hps_io_gpio_inst_GPIO48
			hps_io_gpio_inst_GPIO53  => hps_0_hps_io_hps_io_gpio_inst_GPIO53,          --                  .hps_io_gpio_inst_GPIO53
			hps_io_gpio_inst_GPIO54  => hps_0_hps_io_hps_io_gpio_inst_GPIO54,          --                  .hps_io_gpio_inst_GPIO54
			hps_io_gpio_inst_GPIO61  => hps_0_hps_io_hps_io_gpio_inst_GPIO61,          --                  .hps_io_gpio_inst_GPIO61
			h2f_rst_n                => hps_0_h2f_reset_reset,                         --         h2f_reset.reset_n
			h2f_axi_clk              => clk_clk,                                       --     h2f_axi_clock.clk
			h2f_AWID                 => hps_0_h2f_axi_master_awid,                     --    h2f_axi_master.awid
			h2f_AWADDR               => hps_0_h2f_axi_master_awaddr,                   --                  .awaddr
			h2f_AWLEN                => hps_0_h2f_axi_master_awlen,                    --                  .awlen
			h2f_AWSIZE               => hps_0_h2f_axi_master_awsize,                   --                  .awsize
			h2f_AWBURST              => hps_0_h2f_axi_master_awburst,                  --                  .awburst
			h2f_AWLOCK               => hps_0_h2f_axi_master_awlock,                   --                  .awlock
			h2f_AWCACHE              => hps_0_h2f_axi_master_awcache,                  --                  .awcache
			h2f_AWPROT               => hps_0_h2f_axi_master_awprot,                   --                  .awprot
			h2f_AWVALID              => hps_0_h2f_axi_master_awvalid,                  --                  .awvalid
			h2f_AWREADY              => hps_0_h2f_axi_master_awready,                  --                  .awready
			h2f_WID                  => hps_0_h2f_axi_master_wid,                      --                  .wid
			h2f_WDATA                => hps_0_h2f_axi_master_wdata,                    --                  .wdata
			h2f_WSTRB                => hps_0_h2f_axi_master_wstrb,                    --                  .wstrb
			h2f_WLAST                => hps_0_h2f_axi_master_wlast,                    --                  .wlast
			h2f_WVALID               => hps_0_h2f_axi_master_wvalid,                   --                  .wvalid
			h2f_WREADY               => hps_0_h2f_axi_master_wready,                   --                  .wready
			h2f_BID                  => hps_0_h2f_axi_master_bid,                      --                  .bid
			h2f_BRESP                => hps_0_h2f_axi_master_bresp,                    --                  .bresp
			h2f_BVALID               => hps_0_h2f_axi_master_bvalid,                   --                  .bvalid
			h2f_BREADY               => hps_0_h2f_axi_master_bready,                   --                  .bready
			h2f_ARID                 => hps_0_h2f_axi_master_arid,                     --                  .arid
			h2f_ARADDR               => hps_0_h2f_axi_master_araddr,                   --                  .araddr
			h2f_ARLEN                => hps_0_h2f_axi_master_arlen,                    --                  .arlen
			h2f_ARSIZE               => hps_0_h2f_axi_master_arsize,                   --                  .arsize
			h2f_ARBURST              => hps_0_h2f_axi_master_arburst,                  --                  .arburst
			h2f_ARLOCK               => hps_0_h2f_axi_master_arlock,                   --                  .arlock
			h2f_ARCACHE              => hps_0_h2f_axi_master_arcache,                  --                  .arcache
			h2f_ARPROT               => hps_0_h2f_axi_master_arprot,                   --                  .arprot
			h2f_ARVALID              => hps_0_h2f_axi_master_arvalid,                  --                  .arvalid
			h2f_ARREADY              => hps_0_h2f_axi_master_arready,                  --                  .arready
			h2f_RID                  => hps_0_h2f_axi_master_rid,                      --                  .rid
			h2f_RDATA                => hps_0_h2f_axi_master_rdata,                    --                  .rdata
			h2f_RRESP                => hps_0_h2f_axi_master_rresp,                    --                  .rresp
			h2f_RLAST                => hps_0_h2f_axi_master_rlast,                    --                  .rlast
			h2f_RVALID               => hps_0_h2f_axi_master_rvalid,                   --                  .rvalid
			h2f_RREADY               => hps_0_h2f_axi_master_rready,                   --                  .rready
			f2h_axi_clk              => clk_clk,                                       --     f2h_axi_clock.clk
			f2h_AWID                 => mm_interconnect_0_hps_0_f2h_axi_slave_awid,    --     f2h_axi_slave.awid
			f2h_AWADDR               => mm_interconnect_0_hps_0_f2h_axi_slave_awaddr,  --                  .awaddr
			f2h_AWLEN                => mm_interconnect_0_hps_0_f2h_axi_slave_awlen,   --                  .awlen
			f2h_AWSIZE               => mm_interconnect_0_hps_0_f2h_axi_slave_awsize,  --                  .awsize
			f2h_AWBURST              => mm_interconnect_0_hps_0_f2h_axi_slave_awburst, --                  .awburst
			f2h_AWLOCK               => mm_interconnect_0_hps_0_f2h_axi_slave_awlock,  --                  .awlock
			f2h_AWCACHE              => mm_interconnect_0_hps_0_f2h_axi_slave_awcache, --                  .awcache
			f2h_AWPROT               => mm_interconnect_0_hps_0_f2h_axi_slave_awprot,  --                  .awprot
			f2h_AWVALID              => mm_interconnect_0_hps_0_f2h_axi_slave_awvalid, --                  .awvalid
			f2h_AWREADY              => mm_interconnect_0_hps_0_f2h_axi_slave_awready, --                  .awready
			f2h_AWUSER               => mm_interconnect_0_hps_0_f2h_axi_slave_awuser,  --                  .awuser
			f2h_WID                  => mm_interconnect_0_hps_0_f2h_axi_slave_wid,     --                  .wid
			f2h_WDATA                => mm_interconnect_0_hps_0_f2h_axi_slave_wdata,   --                  .wdata
			f2h_WSTRB                => mm_interconnect_0_hps_0_f2h_axi_slave_wstrb,   --                  .wstrb
			f2h_WLAST                => mm_interconnect_0_hps_0_f2h_axi_slave_wlast,   --                  .wlast
			f2h_WVALID               => mm_interconnect_0_hps_0_f2h_axi_slave_wvalid,  --                  .wvalid
			f2h_WREADY               => mm_interconnect_0_hps_0_f2h_axi_slave_wready,  --                  .wready
			f2h_BID                  => mm_interconnect_0_hps_0_f2h_axi_slave_bid,     --                  .bid
			f2h_BRESP                => mm_interconnect_0_hps_0_f2h_axi_slave_bresp,   --                  .bresp
			f2h_BVALID               => mm_interconnect_0_hps_0_f2h_axi_slave_bvalid,  --                  .bvalid
			f2h_BREADY               => mm_interconnect_0_hps_0_f2h_axi_slave_bready,  --                  .bready
			f2h_ARID                 => mm_interconnect_0_hps_0_f2h_axi_slave_arid,    --                  .arid
			f2h_ARADDR               => mm_interconnect_0_hps_0_f2h_axi_slave_araddr,  --                  .araddr
			f2h_ARLEN                => mm_interconnect_0_hps_0_f2h_axi_slave_arlen,   --                  .arlen
			f2h_ARSIZE               => mm_interconnect_0_hps_0_f2h_axi_slave_arsize,  --                  .arsize
			f2h_ARBURST              => mm_interconnect_0_hps_0_f2h_axi_slave_arburst, --                  .arburst
			f2h_ARLOCK               => mm_interconnect_0_hps_0_f2h_axi_slave_arlock,  --                  .arlock
			f2h_ARCACHE              => mm_interconnect_0_hps_0_f2h_axi_slave_arcache, --                  .arcache
			f2h_ARPROT               => mm_interconnect_0_hps_0_f2h_axi_slave_arprot,  --                  .arprot
			f2h_ARVALID              => mm_interconnect_0_hps_0_f2h_axi_slave_arvalid, --                  .arvalid
			f2h_ARREADY              => mm_interconnect_0_hps_0_f2h_axi_slave_arready, --                  .arready
			f2h_ARUSER               => mm_interconnect_0_hps_0_f2h_axi_slave_aruser,  --                  .aruser
			f2h_RID                  => mm_interconnect_0_hps_0_f2h_axi_slave_rid,     --                  .rid
			f2h_RDATA                => mm_interconnect_0_hps_0_f2h_axi_slave_rdata,   --                  .rdata
			f2h_RRESP                => mm_interconnect_0_hps_0_f2h_axi_slave_rresp,   --                  .rresp
			f2h_RLAST                => mm_interconnect_0_hps_0_f2h_axi_slave_rlast,   --                  .rlast
			f2h_RVALID               => mm_interconnect_0_hps_0_f2h_axi_slave_rvalid,  --                  .rvalid
			f2h_RREADY               => mm_interconnect_0_hps_0_f2h_axi_slave_rready,  --                  .rready
			h2f_lw_axi_clk           => clk_clk,                                       --  h2f_lw_axi_clock.clk
			h2f_lw_AWID              => hps_0_h2f_lw_axi_master_awid,                  -- h2f_lw_axi_master.awid
			h2f_lw_AWADDR            => hps_0_h2f_lw_axi_master_awaddr,                --                  .awaddr
			h2f_lw_AWLEN             => hps_0_h2f_lw_axi_master_awlen,                 --                  .awlen
			h2f_lw_AWSIZE            => hps_0_h2f_lw_axi_master_awsize,                --                  .awsize
			h2f_lw_AWBURST           => hps_0_h2f_lw_axi_master_awburst,               --                  .awburst
			h2f_lw_AWLOCK            => hps_0_h2f_lw_axi_master_awlock,                --                  .awlock
			h2f_lw_AWCACHE           => hps_0_h2f_lw_axi_master_awcache,               --                  .awcache
			h2f_lw_AWPROT            => hps_0_h2f_lw_axi_master_awprot,                --                  .awprot
			h2f_lw_AWVALID           => hps_0_h2f_lw_axi_master_awvalid,               --                  .awvalid
			h2f_lw_AWREADY           => hps_0_h2f_lw_axi_master_awready,               --                  .awready
			h2f_lw_WID               => hps_0_h2f_lw_axi_master_wid,                   --                  .wid
			h2f_lw_WDATA             => hps_0_h2f_lw_axi_master_wdata,                 --                  .wdata
			h2f_lw_WSTRB             => hps_0_h2f_lw_axi_master_wstrb,                 --                  .wstrb
			h2f_lw_WLAST             => hps_0_h2f_lw_axi_master_wlast,                 --                  .wlast
			h2f_lw_WVALID            => hps_0_h2f_lw_axi_master_wvalid,                --                  .wvalid
			h2f_lw_WREADY            => hps_0_h2f_lw_axi_master_wready,                --                  .wready
			h2f_lw_BID               => hps_0_h2f_lw_axi_master_bid,                   --                  .bid
			h2f_lw_BRESP             => hps_0_h2f_lw_axi_master_bresp,                 --                  .bresp
			h2f_lw_BVALID            => hps_0_h2f_lw_axi_master_bvalid,                --                  .bvalid
			h2f_lw_BREADY            => hps_0_h2f_lw_axi_master_bready,                --                  .bready
			h2f_lw_ARID              => hps_0_h2f_lw_axi_master_arid,                  --                  .arid
			h2f_lw_ARADDR            => hps_0_h2f_lw_axi_master_araddr,                --                  .araddr
			h2f_lw_ARLEN             => hps_0_h2f_lw_axi_master_arlen,                 --                  .arlen
			h2f_lw_ARSIZE            => hps_0_h2f_lw_axi_master_arsize,                --                  .arsize
			h2f_lw_ARBURST           => hps_0_h2f_lw_axi_master_arburst,               --                  .arburst
			h2f_lw_ARLOCK            => hps_0_h2f_lw_axi_master_arlock,                --                  .arlock
			h2f_lw_ARCACHE           => hps_0_h2f_lw_axi_master_arcache,               --                  .arcache
			h2f_lw_ARPROT            => hps_0_h2f_lw_axi_master_arprot,                --                  .arprot
			h2f_lw_ARVALID           => hps_0_h2f_lw_axi_master_arvalid,               --                  .arvalid
			h2f_lw_ARREADY           => hps_0_h2f_lw_axi_master_arready,               --                  .arready
			h2f_lw_RID               => hps_0_h2f_lw_axi_master_rid,                   --                  .rid
			h2f_lw_RDATA             => hps_0_h2f_lw_axi_master_rdata,                 --                  .rdata
			h2f_lw_RRESP             => hps_0_h2f_lw_axi_master_rresp,                 --                  .rresp
			h2f_lw_RLAST             => hps_0_h2f_lw_axi_master_rlast,                 --                  .rlast
			h2f_lw_RVALID            => hps_0_h2f_lw_axi_master_rvalid,                --                  .rvalid
			h2f_lw_RREADY            => hps_0_h2f_lw_axi_master_rready,                --                  .rready
			f2h_irq_p0               => hps_0_f2h_irq0_irq,                            --          f2h_irq0.irq
			f2h_irq_p1               => hps_0_f2h_irq1_irq                             --          f2h_irq1.irq
		);

	i2c_ext : component altera_avalon_i2c
		generic map (
			USE_AV_ST       => 0,
			FIFO_DEPTH      => 32,
			FIFO_DEPTH_LOG2 => 5
		)
		port map (
			clk       => clk_clk,                                      --            clock.clk
			rst_n     => rst_controller_003_reset_out_reset_ports_inv, --       reset_sink.reset_n
			intr      => irq_mapper_001_receiver1_irq,                 -- interrupt_sender.irq
			addr      => mm_interconnect_1_i2c_ext_csr_address,        --              csr.address
			read      => mm_interconnect_1_i2c_ext_csr_read,           --                 .read
			write     => mm_interconnect_1_i2c_ext_csr_write,          --                 .write
			writedata => mm_interconnect_1_i2c_ext_csr_writedata,      --                 .writedata
			readdata  => mm_interconnect_1_i2c_ext_csr_readdata,       --                 .readdata
			sda_in    => i2c_ext_sda_in,                               --       i2c_serial.sda_in
			scl_in    => i2c_ext_scl_in,                               --                 .scl_in
			sda_oe    => i2c_ext_sda_oe,                               --                 .sda_oe
			scl_oe    => i2c_ext_scl_oe,                               --                 .scl_oe
			src_data  => open,                                         --      (terminated)
			src_valid => open,                                         --      (terminated)
			src_ready => '0',                                          --      (terminated)
			snk_data  => "0000000000000000",                           --      (terminated)
			snk_valid => '0',                                          --      (terminated)
			snk_ready => open                                          --      (terminated)
		);

	i2c_int : component altera_avalon_i2c
		generic map (
			USE_AV_ST       => 0,
			FIFO_DEPTH      => 32,
			FIFO_DEPTH_LOG2 => 5
		)
		port map (
			clk       => clk_clk,                                      --            clock.clk
			rst_n     => rst_controller_003_reset_out_reset_ports_inv, --       reset_sink.reset_n
			intr      => irq_mapper_001_receiver0_irq,                 -- interrupt_sender.irq
			addr      => mm_interconnect_1_i2c_int_csr_address,        --              csr.address
			read      => mm_interconnect_1_i2c_int_csr_read,           --                 .read
			write     => mm_interconnect_1_i2c_int_csr_write,          --                 .write
			writedata => mm_interconnect_1_i2c_int_csr_writedata,      --                 .writedata
			readdata  => mm_interconnect_1_i2c_int_csr_readdata,       --                 .readdata
			sda_in    => i2c_int_sda_in,                               --       i2c_serial.sda_in
			scl_in    => i2c_int_scl_in,                               --                 .scl_in
			sda_oe    => i2c_int_sda_oe,                               --                 .sda_oe
			scl_oe    => i2c_int_scl_oe,                               --                 .scl_oe
			src_data  => open,                                         --      (terminated)
			src_valid => open,                                         --      (terminated)
			src_ready => '0',                                          --      (terminated)
			snk_data  => "0000000000000000",                           --      (terminated)
			snk_valid => '0',                                          --      (terminated)
			snk_ready => open                                          --      (terminated)
		);

	jtag_uart : component soc_system_v5_jtag_uart
		port map (
			clk            => clk_clk,                                                       --               clk.clk
			rst_n          => rst_controller_003_reset_out_reset_ports_inv,                  --             reset.reset_n
			av_chipselect  => mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_1_jtag_uart_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_1_jtag_uart_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_1_jtag_uart_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver1_irq                                       --               irq.irq
		);

	master_non_sec : component soc_system_v5_master_non_sec
		generic map (
			USE_PLI     => 0,
			PLI_PORT    => 50000,
			FIFO_DEPTHS => 2
		)
		port map (
			clk_clk              => clk_clk,                             --          clk.clk
			clk_reset_reset      => reset_reset_n_ports_inv,             --    clk_reset.reset
			master_address       => master_non_sec_master_address,       --       master.address
			master_readdata      => master_non_sec_master_readdata,      --             .readdata
			master_read          => master_non_sec_master_read,          --             .read
			master_write         => master_non_sec_master_write,         --             .write
			master_writedata     => master_non_sec_master_writedata,     --             .writedata
			master_waitrequest   => master_non_sec_master_waitrequest,   --             .waitrequest
			master_readdatavalid => master_non_sec_master_readdatavalid, --             .readdatavalid
			master_byteenable    => master_non_sec_master_byteenable,    --             .byteenable
			master_reset_reset   => open                                 -- master_reset.reset
		);

	master_secure : component soc_system_v5_master_non_sec
		generic map (
			USE_PLI     => 0,
			PLI_PORT    => 50000,
			FIFO_DEPTHS => 2
		)
		port map (
			clk_clk              => clk_clk,                            --          clk.clk
			clk_reset_reset      => reset_reset_n_ports_inv,            --    clk_reset.reset
			master_address       => master_secure_master_address,       --       master.address
			master_readdata      => master_secure_master_readdata,      --             .readdata
			master_read          => master_secure_master_read,          --             .read
			master_write         => master_secure_master_write,         --             .write
			master_writedata     => master_secure_master_writedata,     --             .writedata
			master_waitrequest   => master_secure_master_waitrequest,   --             .waitrequest
			master_readdatavalid => master_secure_master_readdatavalid, --             .readdatavalid
			master_byteenable    => master_secure_master_byteenable,    --             .byteenable
			master_reset_reset   => open                                -- master_reset.reset
		);

	nmr_parameters : component soc_system_v5_nmr_parameters
		port map (
			adc_val_sub_clk_clk                         => clk_clk,                                                              --                      adc_val_sub_clk.clk
			adc_val_sub_external_connection_export      => adc_val_sub_export,                                                   --      adc_val_sub_external_connection.export
			adc_val_sub_reset_reset_n                   => rst_controller_003_reset_out_reset_ports_inv,                         --                    adc_val_sub_reset.reset_n
			adc_val_sub_s1_address                      => mm_interconnect_1_nmr_parameters_adc_val_sub_s1_address,              --                       adc_val_sub_s1.address
			adc_val_sub_s1_write_n                      => mm_interconnect_1_nmr_parameters_adc_val_sub_s1_write_ports_inv,      --                                     .write_n
			adc_val_sub_s1_writedata                    => mm_interconnect_1_nmr_parameters_adc_val_sub_s1_writedata,            --                                     .writedata
			adc_val_sub_s1_chipselect                   => mm_interconnect_1_nmr_parameters_adc_val_sub_s1_chipselect,           --                                     .chipselect
			adc_val_sub_s1_readdata                     => mm_interconnect_1_nmr_parameters_adc_val_sub_s1_readdata,             --                                     .readdata
			delay_nosig_clk_clk                         => clk_clk,                                                              --                      delay_nosig_clk.clk
			delay_nosig_external_connection_export      => delay_nosig_export,                                                   --      delay_nosig_external_connection.export
			delay_nosig_reset_reset_n                   => rst_controller_003_reset_out_reset_ports_inv,                         --                    delay_nosig_reset.reset_n
			delay_nosig_s1_address                      => mm_interconnect_1_nmr_parameters_delay_nosig_s1_address,              --                       delay_nosig_s1.address
			delay_nosig_s1_write_n                      => mm_interconnect_1_nmr_parameters_delay_nosig_s1_write_ports_inv,      --                                     .write_n
			delay_nosig_s1_writedata                    => mm_interconnect_1_nmr_parameters_delay_nosig_s1_writedata,            --                                     .writedata
			delay_nosig_s1_chipselect                   => mm_interconnect_1_nmr_parameters_delay_nosig_s1_chipselect,           --                                     .chipselect
			delay_nosig_s1_readdata                     => mm_interconnect_1_nmr_parameters_delay_nosig_s1_readdata,             --                                     .readdata
			delay_sig_clk_clk                           => clk_clk,                                                              --                        delay_sig_clk.clk
			delay_sig_external_connection_export        => delay_sig_export,                                                     --        delay_sig_external_connection.export
			delay_sig_reset_reset_n                     => rst_controller_003_reset_out_reset_ports_inv,                         --                      delay_sig_reset.reset_n
			delay_sig_s1_address                        => mm_interconnect_1_nmr_parameters_delay_sig_s1_address,                --                         delay_sig_s1.address
			delay_sig_s1_write_n                        => mm_interconnect_1_nmr_parameters_delay_sig_s1_write_ports_inv,        --                                     .write_n
			delay_sig_s1_writedata                      => mm_interconnect_1_nmr_parameters_delay_sig_s1_writedata,              --                                     .writedata
			delay_sig_s1_chipselect                     => mm_interconnect_1_nmr_parameters_delay_sig_s1_chipselect,             --                                     .chipselect
			delay_sig_s1_readdata                       => mm_interconnect_1_nmr_parameters_delay_sig_s1_readdata,               --                                     .readdata
			delay_t1_clk_clk                            => clk_clk,                                                              --                         delay_t1_clk.clk
			delay_t1_external_connection_export         => delay_t1_export,                                                      --         delay_t1_external_connection.export
			delay_t1_reset_reset_n                      => rst_controller_003_reset_out_reset_ports_inv,                         --                       delay_t1_reset.reset_n
			delay_t1_s1_address                         => mm_interconnect_1_nmr_parameters_delay_t1_s1_address,                 --                          delay_t1_s1.address
			delay_t1_s1_write_n                         => mm_interconnect_1_nmr_parameters_delay_t1_s1_write_ports_inv,         --                                     .write_n
			delay_t1_s1_writedata                       => mm_interconnect_1_nmr_parameters_delay_t1_s1_writedata,               --                                     .writedata
			delay_t1_s1_chipselect                      => mm_interconnect_1_nmr_parameters_delay_t1_s1_chipselect,              --                                     .chipselect
			delay_t1_s1_readdata                        => mm_interconnect_1_nmr_parameters_delay_t1_s1_readdata,                --                                     .readdata
			echoes_per_scan_clk_clk                     => clk_clk,                                                              --                  echoes_per_scan_clk.clk
			echoes_per_scan_external_connection_export  => echoes_per_scan_export,                                               --  echoes_per_scan_external_connection.export
			echoes_per_scan_reset_reset_n               => rst_controller_003_reset_out_reset_ports_inv,                         --                echoes_per_scan_reset.reset_n
			echoes_per_scan_s1_address                  => mm_interconnect_1_nmr_parameters_echoes_per_scan_s1_address,          --                   echoes_per_scan_s1.address
			echoes_per_scan_s1_write_n                  => mm_interconnect_1_nmr_parameters_echoes_per_scan_s1_write_ports_inv,  --                                     .write_n
			echoes_per_scan_s1_writedata                => mm_interconnect_1_nmr_parameters_echoes_per_scan_s1_writedata,        --                                     .writedata
			echoes_per_scan_s1_chipselect               => mm_interconnect_1_nmr_parameters_echoes_per_scan_s1_chipselect,       --                                     .chipselect
			echoes_per_scan_s1_readdata                 => mm_interconnect_1_nmr_parameters_echoes_per_scan_s1_readdata,         --                                     .readdata
			init_delay_clk_clk                          => clk_clk,                                                              --                       init_delay_clk.clk
			init_delay_external_connection_export       => init_delay_export,                                                    --       init_delay_external_connection.export
			init_delay_reset_reset_n                    => rst_controller_003_reset_out_reset_ports_inv,                         --                     init_delay_reset.reset_n
			init_delay_s1_address                       => mm_interconnect_1_nmr_parameters_init_delay_s1_address,               --                        init_delay_s1.address
			init_delay_s1_write_n                       => mm_interconnect_1_nmr_parameters_init_delay_s1_write_ports_inv,       --                                     .write_n
			init_delay_s1_writedata                     => mm_interconnect_1_nmr_parameters_init_delay_s1_writedata,             --                                     .writedata
			init_delay_s1_chipselect                    => mm_interconnect_1_nmr_parameters_init_delay_s1_chipselect,            --                                     .chipselect
			init_delay_s1_readdata                      => mm_interconnect_1_nmr_parameters_init_delay_s1_readdata,              --                                     .readdata
			pulse_180deg_clk_clk                        => clk_clk,                                                              --                     pulse_180deg_clk.clk
			pulse_180deg_external_connection_export     => pulse_180deg_export,                                                  --     pulse_180deg_external_connection.export
			pulse_180deg_reset_reset_n                  => rst_controller_003_reset_out_reset_ports_inv,                         --                   pulse_180deg_reset.reset_n
			pulse_180deg_s1_address                     => mm_interconnect_1_nmr_parameters_pulse_180deg_s1_address,             --                      pulse_180deg_s1.address
			pulse_180deg_s1_write_n                     => mm_interconnect_1_nmr_parameters_pulse_180deg_s1_write_ports_inv,     --                                     .write_n
			pulse_180deg_s1_writedata                   => mm_interconnect_1_nmr_parameters_pulse_180deg_s1_writedata,           --                                     .writedata
			pulse_180deg_s1_chipselect                  => mm_interconnect_1_nmr_parameters_pulse_180deg_s1_chipselect,          --                                     .chipselect
			pulse_180deg_s1_readdata                    => mm_interconnect_1_nmr_parameters_pulse_180deg_s1_readdata,            --                                     .readdata
			pulse_90deg_clk_clk                         => clk_clk,                                                              --                      pulse_90deg_clk.clk
			pulse_90deg_external_connection_export      => pulse_90deg_export,                                                   --      pulse_90deg_external_connection.export
			pulse_90deg_reset_reset_n                   => rst_controller_003_reset_out_reset_ports_inv,                         --                    pulse_90deg_reset.reset_n
			pulse_90deg_s1_address                      => mm_interconnect_1_nmr_parameters_pulse_90deg_s1_address,              --                       pulse_90deg_s1.address
			pulse_90deg_s1_write_n                      => mm_interconnect_1_nmr_parameters_pulse_90deg_s1_write_ports_inv,      --                                     .write_n
			pulse_90deg_s1_writedata                    => mm_interconnect_1_nmr_parameters_pulse_90deg_s1_writedata,            --                                     .writedata
			pulse_90deg_s1_chipselect                   => mm_interconnect_1_nmr_parameters_pulse_90deg_s1_chipselect,           --                                     .chipselect
			pulse_90deg_s1_readdata                     => mm_interconnect_1_nmr_parameters_pulse_90deg_s1_readdata,             --                                     .readdata
			pulse_t1_clk_clk                            => clk_clk,                                                              --                         pulse_t1_clk.clk
			pulse_t1_external_connection_export         => pulse_t1_export,                                                      --         pulse_t1_external_connection.export
			pulse_t1_reset_reset_n                      => rst_controller_003_reset_out_reset_ports_inv,                         --                       pulse_t1_reset.reset_n
			pulse_t1_s1_address                         => mm_interconnect_1_nmr_parameters_pulse_t1_s1_address,                 --                          pulse_t1_s1.address
			pulse_t1_s1_write_n                         => mm_interconnect_1_nmr_parameters_pulse_t1_s1_write_ports_inv,         --                                     .write_n
			pulse_t1_s1_writedata                       => mm_interconnect_1_nmr_parameters_pulse_t1_s1_writedata,               --                                     .writedata
			pulse_t1_s1_chipselect                      => mm_interconnect_1_nmr_parameters_pulse_t1_s1_chipselect,              --                                     .chipselect
			pulse_t1_s1_readdata                        => mm_interconnect_1_nmr_parameters_pulse_t1_s1_readdata,                --                                     .readdata
			rx_delay_clk_clk                            => clk_clk,                                                              --                         rx_delay_clk.clk
			rx_delay_external_connection_export         => rx_delay_export,                                                      --         rx_delay_external_connection.export
			rx_delay_reset_reset_n                      => rst_controller_003_reset_out_reset_ports_inv,                         --                       rx_delay_reset.reset_n
			rx_delay_s1_address                         => mm_interconnect_1_nmr_parameters_rx_delay_s1_address,                 --                          rx_delay_s1.address
			rx_delay_s1_write_n                         => mm_interconnect_1_nmr_parameters_rx_delay_s1_write_ports_inv,         --                                     .write_n
			rx_delay_s1_writedata                       => mm_interconnect_1_nmr_parameters_rx_delay_s1_writedata,               --                                     .writedata
			rx_delay_s1_chipselect                      => mm_interconnect_1_nmr_parameters_rx_delay_s1_chipselect,              --                                     .chipselect
			rx_delay_s1_readdata                        => mm_interconnect_1_nmr_parameters_rx_delay_s1_readdata,                --                                     .readdata
			samples_per_echo_clk_clk                    => clk_clk,                                                              --                 samples_per_echo_clk.clk
			samples_per_echo_external_connection_export => samples_per_echo_export,                                              -- samples_per_echo_external_connection.export
			samples_per_echo_reset_reset_n              => rst_controller_003_reset_out_reset_ports_inv,                         --               samples_per_echo_reset.reset_n
			samples_per_echo_s1_address                 => mm_interconnect_1_nmr_parameters_samples_per_echo_s1_address,         --                  samples_per_echo_s1.address
			samples_per_echo_s1_write_n                 => mm_interconnect_1_nmr_parameters_samples_per_echo_s1_write_ports_inv, --                                     .write_n
			samples_per_echo_s1_writedata               => mm_interconnect_1_nmr_parameters_samples_per_echo_s1_writedata,       --                                     .writedata
			samples_per_echo_s1_chipselect              => mm_interconnect_1_nmr_parameters_samples_per_echo_s1_chipselect,      --                                     .chipselect
			samples_per_echo_s1_readdata                => mm_interconnect_1_nmr_parameters_samples_per_echo_s1_readdata         --                                     .readdata
		);

	nmr_sys_pll : component soc_system_v5_nmr_sys_pll
		port map (
			refclk            => clk_clk,                                              --            refclk.clk
			rst               => nmr_sys_pll_reset_reset,                              --             reset.reset
			outclk_0          => nmr_sys_pll_outclk_clk,                               --           outclk0.clk
			locked            => nmr_sys_pll_locked_export,                            --            locked.export
			reconfig_to_pll   => nmr_sys_pll_reconfig_reconfig_to_pll_reconfig_to_pll, --   reconfig_to_pll.reconfig_to_pll
			reconfig_from_pll => nmr_sys_pll_reconfig_from_pll_reconfig_from_pll       -- reconfig_from_pll.reconfig_from_pll
		);

	nmr_sys_pll_reconfig : component altera_pll_reconfig_top
		generic map (
			device_family       => "Cyclone V",
			ENABLE_MIF          => false,
			MIF_FILE_NAME       => "",
			ENABLE_BYTEENABLE   => false,
			BYTEENABLE_WIDTH    => 4,
			RECONFIG_ADDR_WIDTH => 6,
			RECONFIG_DATA_WIDTH => 32,
			reconf_width        => 64,
			WAIT_FOR_LOCK       => true
		)
		port map (
			mgmt_clk          => clk_clk,                                                              --          mgmt_clk.clk
			mgmt_reset        => rst_controller_003_reset_out_reset,                                   --        mgmt_reset.reset
			mgmt_waitrequest  => mm_interconnect_1_nmr_sys_pll_reconfig_mgmt_avalon_slave_waitrequest, -- mgmt_avalon_slave.waitrequest
			mgmt_read         => mm_interconnect_1_nmr_sys_pll_reconfig_mgmt_avalon_slave_read,        --                  .read
			mgmt_write        => mm_interconnect_1_nmr_sys_pll_reconfig_mgmt_avalon_slave_write,       --                  .write
			mgmt_readdata     => mm_interconnect_1_nmr_sys_pll_reconfig_mgmt_avalon_slave_readdata,    --                  .readdata
			mgmt_address      => mm_interconnect_1_nmr_sys_pll_reconfig_mgmt_avalon_slave_address,     --                  .address
			mgmt_writedata    => mm_interconnect_1_nmr_sys_pll_reconfig_mgmt_avalon_slave_writedata,   --                  .writedata
			reconfig_to_pll   => nmr_sys_pll_reconfig_reconfig_to_pll_reconfig_to_pll,                 --   reconfig_to_pll.reconfig_to_pll
			reconfig_from_pll => nmr_sys_pll_reconfig_from_pll_reconfig_from_pll,                      -- reconfig_from_pll.reconfig_from_pll
			mgmt_byteenable   => "0000"                                                                --       (terminated)
		);

	sdram : component soc_system_v5_sdram
		port map (
			clk            => clk_clk,                                         --   clk.clk
			reset_n        => rst_controller_003_reset_out_reset_ports_inv,    -- reset.reset_n
			az_addr        => mm_interconnect_1_sdram_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_1_sdram_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_1_sdram_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_1_sdram_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_1_sdram_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_1_sdram_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_1_sdram_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_1_sdram_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_1_sdram_s1_waitrequest,          --      .waitrequest
			zs_addr        => sdram_wire_addr,                                 --  wire.export
			zs_ba          => sdram_wire_ba,                                   --      .export
			zs_cas_n       => sdram_wire_cas_n,                                --      .export
			zs_cke         => sdram_wire_cke,                                  --      .export
			zs_cs_n        => sdram_wire_cs_n,                                 --      .export
			zs_dq          => sdram_wire_dq,                                   --      .export
			zs_dqm         => sdram_wire_dqm,                                  --      .export
			zs_ras_n       => sdram_wire_ras_n,                                --      .export
			zs_we_n        => sdram_wire_we_n                                  --      .export
		);

	spi_afe_relays : component soc_system_v5_spi_afe_relays
		port map (
			clk           => clk_clk,                                                           --              clk.clk
			reset_n       => rst_controller_003_reset_out_reset_ports_inv,                      --            reset.reset_n
			data_from_cpu => mm_interconnect_1_spi_afe_relays_spi_control_port_writedata,       -- spi_control_port.writedata
			data_to_cpu   => mm_interconnect_1_spi_afe_relays_spi_control_port_readdata,        --                 .readdata
			mem_addr      => mm_interconnect_1_spi_afe_relays_spi_control_port_address,         --                 .address
			read_n        => mm_interconnect_1_spi_afe_relays_spi_control_port_read_ports_inv,  --                 .read_n
			spi_select    => mm_interconnect_1_spi_afe_relays_spi_control_port_chipselect,      --                 .chipselect
			write_n       => mm_interconnect_1_spi_afe_relays_spi_control_port_write_ports_inv, --                 .write_n
			irq           => irq_mapper_001_receiver7_irq,                                      --              irq.irq
			MISO          => spi_afe_relays_MISO,                                               --         external.export
			MOSI          => spi_afe_relays_MOSI,                                               --                 .export
			SCLK          => spi_afe_relays_SCLK,                                               --                 .export
			SS_n          => spi_afe_relays_SS_n                                                --                 .export
		);

	spi_mtch_ntwrk : component soc_system_v5_spi_afe_relays
		port map (
			clk           => clk_clk,                                                           --              clk.clk
			reset_n       => rst_controller_003_reset_out_reset_ports_inv,                      --            reset.reset_n
			data_from_cpu => mm_interconnect_1_spi_mtch_ntwrk_spi_control_port_writedata,       -- spi_control_port.writedata
			data_to_cpu   => mm_interconnect_1_spi_mtch_ntwrk_spi_control_port_readdata,        --                 .readdata
			mem_addr      => mm_interconnect_1_spi_mtch_ntwrk_spi_control_port_address,         --                 .address
			read_n        => mm_interconnect_1_spi_mtch_ntwrk_spi_control_port_read_ports_inv,  --                 .read_n
			spi_select    => mm_interconnect_1_spi_mtch_ntwrk_spi_control_port_chipselect,      --                 .chipselect
			write_n       => mm_interconnect_1_spi_mtch_ntwrk_spi_control_port_write_ports_inv, --                 .write_n
			irq           => irq_mapper_001_receiver4_irq,                                      --              irq.irq
			MISO          => spi_mtch_ntwrk_MISO,                                               --         external.export
			MOSI          => spi_mtch_ntwrk_MOSI,                                               --                 .export
			SCLK          => spi_mtch_ntwrk_SCLK,                                               --                 .export
			SS_n          => spi_mtch_ntwrk_SS_n                                                --                 .export
		);

	switches : component soc_system_v5_switches
		port map (
			clk      => clk_clk,                                      --                 clk.clk
			reset_n  => rst_controller_003_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_1_switches_s1_address,        --                  s1.address
			readdata => mm_interconnect_1_switches_s1_readdata,       --                    .readdata
			in_port  => switches_export                               -- external_connection.export
		);

	sysid_qsys : component soc_system_v5_sysid_qsys
		port map (
			clock    => clk_clk,                                               --           clk.clk
			reset_n  => rst_controller_003_reset_out_reset_ports_inv,          --         reset.reset_n
			readdata => mm_interconnect_1_sysid_qsys_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_1_sysid_qsys_control_slave_address(0)  --              .address
		);

	mm_interconnect_0 : component soc_system_v5_mm_interconnect_0
		port map (
			hps_0_f2h_axi_slave_awid                                         => mm_interconnect_0_hps_0_f2h_axi_slave_awid,    --                                        hps_0_f2h_axi_slave.awid
			hps_0_f2h_axi_slave_awaddr                                       => mm_interconnect_0_hps_0_f2h_axi_slave_awaddr,  --                                                           .awaddr
			hps_0_f2h_axi_slave_awlen                                        => mm_interconnect_0_hps_0_f2h_axi_slave_awlen,   --                                                           .awlen
			hps_0_f2h_axi_slave_awsize                                       => mm_interconnect_0_hps_0_f2h_axi_slave_awsize,  --                                                           .awsize
			hps_0_f2h_axi_slave_awburst                                      => mm_interconnect_0_hps_0_f2h_axi_slave_awburst, --                                                           .awburst
			hps_0_f2h_axi_slave_awlock                                       => mm_interconnect_0_hps_0_f2h_axi_slave_awlock,  --                                                           .awlock
			hps_0_f2h_axi_slave_awcache                                      => mm_interconnect_0_hps_0_f2h_axi_slave_awcache, --                                                           .awcache
			hps_0_f2h_axi_slave_awprot                                       => mm_interconnect_0_hps_0_f2h_axi_slave_awprot,  --                                                           .awprot
			hps_0_f2h_axi_slave_awuser                                       => mm_interconnect_0_hps_0_f2h_axi_slave_awuser,  --                                                           .awuser
			hps_0_f2h_axi_slave_awvalid                                      => mm_interconnect_0_hps_0_f2h_axi_slave_awvalid, --                                                           .awvalid
			hps_0_f2h_axi_slave_awready                                      => mm_interconnect_0_hps_0_f2h_axi_slave_awready, --                                                           .awready
			hps_0_f2h_axi_slave_wid                                          => mm_interconnect_0_hps_0_f2h_axi_slave_wid,     --                                                           .wid
			hps_0_f2h_axi_slave_wdata                                        => mm_interconnect_0_hps_0_f2h_axi_slave_wdata,   --                                                           .wdata
			hps_0_f2h_axi_slave_wstrb                                        => mm_interconnect_0_hps_0_f2h_axi_slave_wstrb,   --                                                           .wstrb
			hps_0_f2h_axi_slave_wlast                                        => mm_interconnect_0_hps_0_f2h_axi_slave_wlast,   --                                                           .wlast
			hps_0_f2h_axi_slave_wvalid                                       => mm_interconnect_0_hps_0_f2h_axi_slave_wvalid,  --                                                           .wvalid
			hps_0_f2h_axi_slave_wready                                       => mm_interconnect_0_hps_0_f2h_axi_slave_wready,  --                                                           .wready
			hps_0_f2h_axi_slave_bid                                          => mm_interconnect_0_hps_0_f2h_axi_slave_bid,     --                                                           .bid
			hps_0_f2h_axi_slave_bresp                                        => mm_interconnect_0_hps_0_f2h_axi_slave_bresp,   --                                                           .bresp
			hps_0_f2h_axi_slave_bvalid                                       => mm_interconnect_0_hps_0_f2h_axi_slave_bvalid,  --                                                           .bvalid
			hps_0_f2h_axi_slave_bready                                       => mm_interconnect_0_hps_0_f2h_axi_slave_bready,  --                                                           .bready
			hps_0_f2h_axi_slave_arid                                         => mm_interconnect_0_hps_0_f2h_axi_slave_arid,    --                                                           .arid
			hps_0_f2h_axi_slave_araddr                                       => mm_interconnect_0_hps_0_f2h_axi_slave_araddr,  --                                                           .araddr
			hps_0_f2h_axi_slave_arlen                                        => mm_interconnect_0_hps_0_f2h_axi_slave_arlen,   --                                                           .arlen
			hps_0_f2h_axi_slave_arsize                                       => mm_interconnect_0_hps_0_f2h_axi_slave_arsize,  --                                                           .arsize
			hps_0_f2h_axi_slave_arburst                                      => mm_interconnect_0_hps_0_f2h_axi_slave_arburst, --                                                           .arburst
			hps_0_f2h_axi_slave_arlock                                       => mm_interconnect_0_hps_0_f2h_axi_slave_arlock,  --                                                           .arlock
			hps_0_f2h_axi_slave_arcache                                      => mm_interconnect_0_hps_0_f2h_axi_slave_arcache, --                                                           .arcache
			hps_0_f2h_axi_slave_arprot                                       => mm_interconnect_0_hps_0_f2h_axi_slave_arprot,  --                                                           .arprot
			hps_0_f2h_axi_slave_aruser                                       => mm_interconnect_0_hps_0_f2h_axi_slave_aruser,  --                                                           .aruser
			hps_0_f2h_axi_slave_arvalid                                      => mm_interconnect_0_hps_0_f2h_axi_slave_arvalid, --                                                           .arvalid
			hps_0_f2h_axi_slave_arready                                      => mm_interconnect_0_hps_0_f2h_axi_slave_arready, --                                                           .arready
			hps_0_f2h_axi_slave_rid                                          => mm_interconnect_0_hps_0_f2h_axi_slave_rid,     --                                                           .rid
			hps_0_f2h_axi_slave_rdata                                        => mm_interconnect_0_hps_0_f2h_axi_slave_rdata,   --                                                           .rdata
			hps_0_f2h_axi_slave_rresp                                        => mm_interconnect_0_hps_0_f2h_axi_slave_rresp,   --                                                           .rresp
			hps_0_f2h_axi_slave_rlast                                        => mm_interconnect_0_hps_0_f2h_axi_slave_rlast,   --                                                           .rlast
			hps_0_f2h_axi_slave_rvalid                                       => mm_interconnect_0_hps_0_f2h_axi_slave_rvalid,  --                                                           .rvalid
			hps_0_f2h_axi_slave_rready                                       => mm_interconnect_0_hps_0_f2h_axi_slave_rready,  --                                                           .rready
			clk_0_clk_clk                                                    => clk_clk,                                       --                                                  clk_0_clk.clk
			alt_vip_vfr_vga_clock_master_reset_reset_bridge_in_reset_reset   => rst_controller_003_reset_out_reset,            --   alt_vip_vfr_vga_clock_master_reset_reset_bridge_in_reset.reset
			hps_0_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset_reset => rst_controller_004_reset_out_reset,            -- hps_0_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset.reset
			master_secure_clk_reset_reset_bridge_in_reset_reset              => rst_controller_003_reset_out_reset,            --              master_secure_clk_reset_reset_bridge_in_reset.reset
			alt_vip_vfr_vga_avalon_master_address                            => alt_vip_vfr_vga_avalon_master_address,         --                              alt_vip_vfr_vga_avalon_master.address
			alt_vip_vfr_vga_avalon_master_waitrequest                        => alt_vip_vfr_vga_avalon_master_waitrequest,     --                                                           .waitrequest
			alt_vip_vfr_vga_avalon_master_burstcount                         => alt_vip_vfr_vga_avalon_master_burstcount,      --                                                           .burstcount
			alt_vip_vfr_vga_avalon_master_read                               => alt_vip_vfr_vga_avalon_master_read,            --                                                           .read
			alt_vip_vfr_vga_avalon_master_readdata                           => alt_vip_vfr_vga_avalon_master_readdata,        --                                                           .readdata
			alt_vip_vfr_vga_avalon_master_readdatavalid                      => alt_vip_vfr_vga_avalon_master_readdatavalid,   --                                                           .readdatavalid
			master_secure_master_address                                     => master_secure_master_address,                  --                                       master_secure_master.address
			master_secure_master_waitrequest                                 => master_secure_master_waitrequest,              --                                                           .waitrequest
			master_secure_master_byteenable                                  => master_secure_master_byteenable,               --                                                           .byteenable
			master_secure_master_read                                        => master_secure_master_read,                     --                                                           .read
			master_secure_master_readdata                                    => master_secure_master_readdata,                 --                                                           .readdata
			master_secure_master_readdatavalid                               => master_secure_master_readdatavalid,            --                                                           .readdatavalid
			master_secure_master_write                                       => master_secure_master_write,                    --                                                           .write
			master_secure_master_writedata                                   => master_secure_master_writedata                 --                                                           .writedata
		);

	mm_interconnect_1 : component soc_system_v5_mm_interconnect_1
		port map (
			hps_0_h2f_axi_master_awid                                        => hps_0_h2f_axi_master_awid,                                             --                                       hps_0_h2f_axi_master.awid
			hps_0_h2f_axi_master_awaddr                                      => hps_0_h2f_axi_master_awaddr,                                           --                                                           .awaddr
			hps_0_h2f_axi_master_awlen                                       => hps_0_h2f_axi_master_awlen,                                            --                                                           .awlen
			hps_0_h2f_axi_master_awsize                                      => hps_0_h2f_axi_master_awsize,                                           --                                                           .awsize
			hps_0_h2f_axi_master_awburst                                     => hps_0_h2f_axi_master_awburst,                                          --                                                           .awburst
			hps_0_h2f_axi_master_awlock                                      => hps_0_h2f_axi_master_awlock,                                           --                                                           .awlock
			hps_0_h2f_axi_master_awcache                                     => hps_0_h2f_axi_master_awcache,                                          --                                                           .awcache
			hps_0_h2f_axi_master_awprot                                      => hps_0_h2f_axi_master_awprot,                                           --                                                           .awprot
			hps_0_h2f_axi_master_awvalid                                     => hps_0_h2f_axi_master_awvalid,                                          --                                                           .awvalid
			hps_0_h2f_axi_master_awready                                     => hps_0_h2f_axi_master_awready,                                          --                                                           .awready
			hps_0_h2f_axi_master_wid                                         => hps_0_h2f_axi_master_wid,                                              --                                                           .wid
			hps_0_h2f_axi_master_wdata                                       => hps_0_h2f_axi_master_wdata,                                            --                                                           .wdata
			hps_0_h2f_axi_master_wstrb                                       => hps_0_h2f_axi_master_wstrb,                                            --                                                           .wstrb
			hps_0_h2f_axi_master_wlast                                       => hps_0_h2f_axi_master_wlast,                                            --                                                           .wlast
			hps_0_h2f_axi_master_wvalid                                      => hps_0_h2f_axi_master_wvalid,                                           --                                                           .wvalid
			hps_0_h2f_axi_master_wready                                      => hps_0_h2f_axi_master_wready,                                           --                                                           .wready
			hps_0_h2f_axi_master_bid                                         => hps_0_h2f_axi_master_bid,                                              --                                                           .bid
			hps_0_h2f_axi_master_bresp                                       => hps_0_h2f_axi_master_bresp,                                            --                                                           .bresp
			hps_0_h2f_axi_master_bvalid                                      => hps_0_h2f_axi_master_bvalid,                                           --                                                           .bvalid
			hps_0_h2f_axi_master_bready                                      => hps_0_h2f_axi_master_bready,                                           --                                                           .bready
			hps_0_h2f_axi_master_arid                                        => hps_0_h2f_axi_master_arid,                                             --                                                           .arid
			hps_0_h2f_axi_master_araddr                                      => hps_0_h2f_axi_master_araddr,                                           --                                                           .araddr
			hps_0_h2f_axi_master_arlen                                       => hps_0_h2f_axi_master_arlen,                                            --                                                           .arlen
			hps_0_h2f_axi_master_arsize                                      => hps_0_h2f_axi_master_arsize,                                           --                                                           .arsize
			hps_0_h2f_axi_master_arburst                                     => hps_0_h2f_axi_master_arburst,                                          --                                                           .arburst
			hps_0_h2f_axi_master_arlock                                      => hps_0_h2f_axi_master_arlock,                                           --                                                           .arlock
			hps_0_h2f_axi_master_arcache                                     => hps_0_h2f_axi_master_arcache,                                          --                                                           .arcache
			hps_0_h2f_axi_master_arprot                                      => hps_0_h2f_axi_master_arprot,                                           --                                                           .arprot
			hps_0_h2f_axi_master_arvalid                                     => hps_0_h2f_axi_master_arvalid,                                          --                                                           .arvalid
			hps_0_h2f_axi_master_arready                                     => hps_0_h2f_axi_master_arready,                                          --                                                           .arready
			hps_0_h2f_axi_master_rid                                         => hps_0_h2f_axi_master_rid,                                              --                                                           .rid
			hps_0_h2f_axi_master_rdata                                       => hps_0_h2f_axi_master_rdata,                                            --                                                           .rdata
			hps_0_h2f_axi_master_rresp                                       => hps_0_h2f_axi_master_rresp,                                            --                                                           .rresp
			hps_0_h2f_axi_master_rlast                                       => hps_0_h2f_axi_master_rlast,                                            --                                                           .rlast
			hps_0_h2f_axi_master_rvalid                                      => hps_0_h2f_axi_master_rvalid,                                           --                                                           .rvalid
			hps_0_h2f_axi_master_rready                                      => hps_0_h2f_axi_master_rready,                                           --                                                           .rready
			hps_0_h2f_lw_axi_master_awid                                     => hps_0_h2f_lw_axi_master_awid,                                          --                                    hps_0_h2f_lw_axi_master.awid
			hps_0_h2f_lw_axi_master_awaddr                                   => hps_0_h2f_lw_axi_master_awaddr,                                        --                                                           .awaddr
			hps_0_h2f_lw_axi_master_awlen                                    => hps_0_h2f_lw_axi_master_awlen,                                         --                                                           .awlen
			hps_0_h2f_lw_axi_master_awsize                                   => hps_0_h2f_lw_axi_master_awsize,                                        --                                                           .awsize
			hps_0_h2f_lw_axi_master_awburst                                  => hps_0_h2f_lw_axi_master_awburst,                                       --                                                           .awburst
			hps_0_h2f_lw_axi_master_awlock                                   => hps_0_h2f_lw_axi_master_awlock,                                        --                                                           .awlock
			hps_0_h2f_lw_axi_master_awcache                                  => hps_0_h2f_lw_axi_master_awcache,                                       --                                                           .awcache
			hps_0_h2f_lw_axi_master_awprot                                   => hps_0_h2f_lw_axi_master_awprot,                                        --                                                           .awprot
			hps_0_h2f_lw_axi_master_awvalid                                  => hps_0_h2f_lw_axi_master_awvalid,                                       --                                                           .awvalid
			hps_0_h2f_lw_axi_master_awready                                  => hps_0_h2f_lw_axi_master_awready,                                       --                                                           .awready
			hps_0_h2f_lw_axi_master_wid                                      => hps_0_h2f_lw_axi_master_wid,                                           --                                                           .wid
			hps_0_h2f_lw_axi_master_wdata                                    => hps_0_h2f_lw_axi_master_wdata,                                         --                                                           .wdata
			hps_0_h2f_lw_axi_master_wstrb                                    => hps_0_h2f_lw_axi_master_wstrb,                                         --                                                           .wstrb
			hps_0_h2f_lw_axi_master_wlast                                    => hps_0_h2f_lw_axi_master_wlast,                                         --                                                           .wlast
			hps_0_h2f_lw_axi_master_wvalid                                   => hps_0_h2f_lw_axi_master_wvalid,                                        --                                                           .wvalid
			hps_0_h2f_lw_axi_master_wready                                   => hps_0_h2f_lw_axi_master_wready,                                        --                                                           .wready
			hps_0_h2f_lw_axi_master_bid                                      => hps_0_h2f_lw_axi_master_bid,                                           --                                                           .bid
			hps_0_h2f_lw_axi_master_bresp                                    => hps_0_h2f_lw_axi_master_bresp,                                         --                                                           .bresp
			hps_0_h2f_lw_axi_master_bvalid                                   => hps_0_h2f_lw_axi_master_bvalid,                                        --                                                           .bvalid
			hps_0_h2f_lw_axi_master_bready                                   => hps_0_h2f_lw_axi_master_bready,                                        --                                                           .bready
			hps_0_h2f_lw_axi_master_arid                                     => hps_0_h2f_lw_axi_master_arid,                                          --                                                           .arid
			hps_0_h2f_lw_axi_master_araddr                                   => hps_0_h2f_lw_axi_master_araddr,                                        --                                                           .araddr
			hps_0_h2f_lw_axi_master_arlen                                    => hps_0_h2f_lw_axi_master_arlen,                                         --                                                           .arlen
			hps_0_h2f_lw_axi_master_arsize                                   => hps_0_h2f_lw_axi_master_arsize,                                        --                                                           .arsize
			hps_0_h2f_lw_axi_master_arburst                                  => hps_0_h2f_lw_axi_master_arburst,                                       --                                                           .arburst
			hps_0_h2f_lw_axi_master_arlock                                   => hps_0_h2f_lw_axi_master_arlock,                                        --                                                           .arlock
			hps_0_h2f_lw_axi_master_arcache                                  => hps_0_h2f_lw_axi_master_arcache,                                       --                                                           .arcache
			hps_0_h2f_lw_axi_master_arprot                                   => hps_0_h2f_lw_axi_master_arprot,                                        --                                                           .arprot
			hps_0_h2f_lw_axi_master_arvalid                                  => hps_0_h2f_lw_axi_master_arvalid,                                       --                                                           .arvalid
			hps_0_h2f_lw_axi_master_arready                                  => hps_0_h2f_lw_axi_master_arready,                                       --                                                           .arready
			hps_0_h2f_lw_axi_master_rid                                      => hps_0_h2f_lw_axi_master_rid,                                           --                                                           .rid
			hps_0_h2f_lw_axi_master_rdata                                    => hps_0_h2f_lw_axi_master_rdata,                                         --                                                           .rdata
			hps_0_h2f_lw_axi_master_rresp                                    => hps_0_h2f_lw_axi_master_rresp,                                         --                                                           .rresp
			hps_0_h2f_lw_axi_master_rlast                                    => hps_0_h2f_lw_axi_master_rlast,                                         --                                                           .rlast
			hps_0_h2f_lw_axi_master_rvalid                                   => hps_0_h2f_lw_axi_master_rvalid,                                        --                                                           .rvalid
			hps_0_h2f_lw_axi_master_rready                                   => hps_0_h2f_lw_axi_master_rready,                                        --                                                           .rready
			clk_0_clk_clk                                                    => clk_clk,                                                               --                                                  clk_0_clk.clk
			gp_pll_outclk0_clk                                               => gp_pll_outclk0_clk,                                                    --                                             gp_pll_outclk0.clk
			adc_fifo_mem_reset_in_reset_bridge_in_reset_reset                => rst_controller_001_reset_out_reset,                                    --                adc_fifo_mem_reset_in_reset_bridge_in_reset.reset
			alt_vip_vfr_vga_clock_reset_reset_reset_bridge_in_reset_reset    => rst_controller_002_reset_out_reset,                                    --    alt_vip_vfr_vga_clock_reset_reset_reset_bridge_in_reset.reset
			dma_fifo_reset_reset_bridge_in_reset_reset                       => rst_controller_003_reset_out_reset,                                    --                       dma_fifo_reset_reset_bridge_in_reset.reset
			hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset => rst_controller_004_reset_out_reset,                                    -- hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
			master_non_sec_clk_reset_reset_bridge_in_reset_reset             => rst_controller_003_reset_out_reset,                                    --             master_non_sec_clk_reset_reset_bridge_in_reset.reset
			dma_dconvi_read_master_address                                   => dma_dconvi_read_master_address,                                        --                                     dma_dconvi_read_master.address
			dma_dconvi_read_master_waitrequest                               => dma_dconvi_read_master_waitrequest,                                    --                                                           .waitrequest
			dma_dconvi_read_master_chipselect                                => dma_dconvi_read_master_chipselect,                                     --                                                           .chipselect
			dma_dconvi_read_master_read                                      => dma_dconvi_read_master_read_ports_inv,                                 --                                                           .read
			dma_dconvi_read_master_readdata                                  => dma_dconvi_read_master_readdata,                                       --                                                           .readdata
			dma_dconvi_read_master_readdatavalid                             => dma_dconvi_read_master_readdatavalid,                                  --                                                           .readdatavalid
			dma_dconvi_write_master_address                                  => dma_dconvi_write_master_address,                                       --                                    dma_dconvi_write_master.address
			dma_dconvi_write_master_waitrequest                              => dma_dconvi_write_master_waitrequest,                                   --                                                           .waitrequest
			dma_dconvi_write_master_byteenable                               => dma_dconvi_write_master_byteenable,                                    --                                                           .byteenable
			dma_dconvi_write_master_chipselect                               => dma_dconvi_write_master_chipselect,                                    --                                                           .chipselect
			dma_dconvi_write_master_write                                    => dma_dconvi_write_master_write_ports_inv,                               --                                                           .write
			dma_dconvi_write_master_writedata                                => dma_dconvi_write_master_writedata,                                     --                                                           .writedata
			dma_dconvq_read_master_address                                   => dma_dconvq_read_master_address,                                        --                                     dma_dconvq_read_master.address
			dma_dconvq_read_master_waitrequest                               => dma_dconvq_read_master_waitrequest,                                    --                                                           .waitrequest
			dma_dconvq_read_master_chipselect                                => dma_dconvq_read_master_chipselect,                                     --                                                           .chipselect
			dma_dconvq_read_master_read                                      => dma_dconvq_read_master_read_ports_inv,                                 --                                                           .read
			dma_dconvq_read_master_readdata                                  => dma_dconvq_read_master_readdata,                                       --                                                           .readdata
			dma_dconvq_read_master_readdatavalid                             => dma_dconvq_read_master_readdatavalid,                                  --                                                           .readdatavalid
			dma_dconvq_write_master_address                                  => dma_dconvq_write_master_address,                                       --                                    dma_dconvq_write_master.address
			dma_dconvq_write_master_waitrequest                              => dma_dconvq_write_master_waitrequest,                                   --                                                           .waitrequest
			dma_dconvq_write_master_byteenable                               => dma_dconvq_write_master_byteenable,                                    --                                                           .byteenable
			dma_dconvq_write_master_chipselect                               => dma_dconvq_write_master_chipselect,                                    --                                                           .chipselect
			dma_dconvq_write_master_write                                    => dma_dconvq_write_master_write_ports_inv,                               --                                                           .write
			dma_dconvq_write_master_writedata                                => dma_dconvq_write_master_writedata,                                     --                                                           .writedata
			dma_dummy_read_master_address                                    => dma_dummy_read_master_address,                                         --                                      dma_dummy_read_master.address
			dma_dummy_read_master_waitrequest                                => dma_dummy_read_master_waitrequest,                                     --                                                           .waitrequest
			dma_dummy_read_master_chipselect                                 => dma_dummy_read_master_chipselect,                                      --                                                           .chipselect
			dma_dummy_read_master_read                                       => dma_dummy_read_master_read_ports_inv,                                  --                                                           .read
			dma_dummy_read_master_readdata                                   => dma_dummy_read_master_readdata,                                        --                                                           .readdata
			dma_dummy_read_master_readdatavalid                              => dma_dummy_read_master_readdatavalid,                                   --                                                           .readdatavalid
			dma_dummy_write_master_address                                   => dma_dummy_write_master_address,                                        --                                     dma_dummy_write_master.address
			dma_dummy_write_master_waitrequest                               => dma_dummy_write_master_waitrequest,                                    --                                                           .waitrequest
			dma_dummy_write_master_byteenable                                => dma_dummy_write_master_byteenable,                                     --                                                           .byteenable
			dma_dummy_write_master_chipselect                                => dma_dummy_write_master_chipselect,                                     --                                                           .chipselect
			dma_dummy_write_master_write                                     => dma_dummy_write_master_write_ports_inv,                                --                                                           .write
			dma_dummy_write_master_writedata                                 => dma_dummy_write_master_writedata,                                      --                                                           .writedata
			dma_fifo_read_master_address                                     => dma_fifo_read_master_address,                                          --                                       dma_fifo_read_master.address
			dma_fifo_read_master_waitrequest                                 => dma_fifo_read_master_waitrequest,                                      --                                                           .waitrequest
			dma_fifo_read_master_chipselect                                  => dma_fifo_read_master_chipselect,                                       --                                                           .chipselect
			dma_fifo_read_master_read                                        => dma_fifo_read_master_read_ports_inv,                                   --                                                           .read
			dma_fifo_read_master_readdata                                    => dma_fifo_read_master_readdata,                                         --                                                           .readdata
			dma_fifo_read_master_readdatavalid                               => dma_fifo_read_master_readdatavalid,                                    --                                                           .readdatavalid
			dma_fifo_write_master_address                                    => dma_fifo_write_master_address,                                         --                                      dma_fifo_write_master.address
			dma_fifo_write_master_waitrequest                                => dma_fifo_write_master_waitrequest,                                     --                                                           .waitrequest
			dma_fifo_write_master_byteenable                                 => dma_fifo_write_master_byteenable,                                      --                                                           .byteenable
			dma_fifo_write_master_chipselect                                 => dma_fifo_write_master_chipselect,                                      --                                                           .chipselect
			dma_fifo_write_master_write                                      => dma_fifo_write_master_write_ports_inv,                                 --                                                           .write
			dma_fifo_write_master_writedata                                  => dma_fifo_write_master_writedata,                                       --                                                           .writedata
			master_non_sec_master_address                                    => master_non_sec_master_address,                                         --                                      master_non_sec_master.address
			master_non_sec_master_waitrequest                                => master_non_sec_master_waitrequest,                                     --                                                           .waitrequest
			master_non_sec_master_byteenable                                 => master_non_sec_master_byteenable,                                      --                                                           .byteenable
			master_non_sec_master_read                                       => master_non_sec_master_read,                                            --                                                           .read
			master_non_sec_master_readdata                                   => master_non_sec_master_readdata,                                        --                                                           .readdata
			master_non_sec_master_readdatavalid                              => master_non_sec_master_readdatavalid,                                   --                                                           .readdatavalid
			master_non_sec_master_write                                      => master_non_sec_master_write,                                           --                                                           .write
			master_non_sec_master_writedata                                  => master_non_sec_master_writedata,                                       --                                                           .writedata
			adc_fifo_mem_in_csr_address                                      => mm_interconnect_1_adc_fifo_mem_in_csr_address,                         --                                        adc_fifo_mem_in_csr.address
			adc_fifo_mem_in_csr_write                                        => mm_interconnect_1_adc_fifo_mem_in_csr_write,                           --                                                           .write
			adc_fifo_mem_in_csr_read                                         => mm_interconnect_1_adc_fifo_mem_in_csr_read,                            --                                                           .read
			adc_fifo_mem_in_csr_readdata                                     => mm_interconnect_1_adc_fifo_mem_in_csr_readdata,                        --                                                           .readdata
			adc_fifo_mem_in_csr_writedata                                    => mm_interconnect_1_adc_fifo_mem_in_csr_writedata,                       --                                                           .writedata
			adc_fifo_mem_out_address                                         => mm_interconnect_1_adc_fifo_mem_out_address,                            --                                           adc_fifo_mem_out.address
			adc_fifo_mem_out_read                                            => mm_interconnect_1_adc_fifo_mem_out_read,                               --                                                           .read
			adc_fifo_mem_out_readdata                                        => mm_interconnect_1_adc_fifo_mem_out_readdata,                           --                                                           .readdata
			adc_fifo_mem_out_waitrequest                                     => mm_interconnect_1_adc_fifo_mem_out_waitrequest,                        --                                                           .waitrequest
			alt_vip_vfr_vga_avalon_slave_address                             => mm_interconnect_1_alt_vip_vfr_vga_avalon_slave_address,                --                               alt_vip_vfr_vga_avalon_slave.address
			alt_vip_vfr_vga_avalon_slave_write                               => mm_interconnect_1_alt_vip_vfr_vga_avalon_slave_write,                  --                                                           .write
			alt_vip_vfr_vga_avalon_slave_read                                => mm_interconnect_1_alt_vip_vfr_vga_avalon_slave_read,                   --                                                           .read
			alt_vip_vfr_vga_avalon_slave_readdata                            => mm_interconnect_1_alt_vip_vfr_vga_avalon_slave_readdata,               --                                                           .readdata
			alt_vip_vfr_vga_avalon_slave_writedata                           => mm_interconnect_1_alt_vip_vfr_vga_avalon_slave_writedata,              --                                                           .writedata
			analyzer_pll_reconfig_mgmt_avalon_slave_address                  => mm_interconnect_1_analyzer_pll_reconfig_mgmt_avalon_slave_address,     --                    analyzer_pll_reconfig_mgmt_avalon_slave.address
			analyzer_pll_reconfig_mgmt_avalon_slave_write                    => mm_interconnect_1_analyzer_pll_reconfig_mgmt_avalon_slave_write,       --                                                           .write
			analyzer_pll_reconfig_mgmt_avalon_slave_read                     => mm_interconnect_1_analyzer_pll_reconfig_mgmt_avalon_slave_read,        --                                                           .read
			analyzer_pll_reconfig_mgmt_avalon_slave_readdata                 => mm_interconnect_1_analyzer_pll_reconfig_mgmt_avalon_slave_readdata,    --                                                           .readdata
			analyzer_pll_reconfig_mgmt_avalon_slave_writedata                => mm_interconnect_1_analyzer_pll_reconfig_mgmt_avalon_slave_writedata,   --                                                           .writedata
			analyzer_pll_reconfig_mgmt_avalon_slave_waitrequest              => mm_interconnect_1_analyzer_pll_reconfig_mgmt_avalon_slave_waitrequest, --                                                           .waitrequest
			aux_cnt_out_s1_address                                           => mm_interconnect_1_aux_cnt_out_s1_address,                              --                                             aux_cnt_out_s1.address
			aux_cnt_out_s1_write                                             => mm_interconnect_1_aux_cnt_out_s1_write,                                --                                                           .write
			aux_cnt_out_s1_readdata                                          => mm_interconnect_1_aux_cnt_out_s1_readdata,                             --                                                           .readdata
			aux_cnt_out_s1_writedata                                         => mm_interconnect_1_aux_cnt_out_s1_writedata,                            --                                                           .writedata
			aux_cnt_out_s1_chipselect                                        => mm_interconnect_1_aux_cnt_out_s1_chipselect,                           --                                                           .chipselect
			ctrl_in_s1_address                                               => mm_interconnect_1_ctrl_in_s1_address,                                  --                                                 ctrl_in_s1.address
			ctrl_in_s1_readdata                                              => mm_interconnect_1_ctrl_in_s1_readdata,                                 --                                                           .readdata
			ctrl_out_s1_address                                              => mm_interconnect_1_ctrl_out_s1_address,                                 --                                                ctrl_out_s1.address
			ctrl_out_s1_write                                                => mm_interconnect_1_ctrl_out_s1_write,                                   --                                                           .write
			ctrl_out_s1_readdata                                             => mm_interconnect_1_ctrl_out_s1_readdata,                                --                                                           .readdata
			ctrl_out_s1_writedata                                            => mm_interconnect_1_ctrl_out_s1_writedata,                               --                                                           .writedata
			ctrl_out_s1_chipselect                                           => mm_interconnect_1_ctrl_out_s1_chipselect,                              --                                                           .chipselect
			dac_grad_spi_control_port_address                                => mm_interconnect_1_dac_grad_spi_control_port_address,                   --                                  dac_grad_spi_control_port.address
			dac_grad_spi_control_port_write                                  => mm_interconnect_1_dac_grad_spi_control_port_write,                     --                                                           .write
			dac_grad_spi_control_port_read                                   => mm_interconnect_1_dac_grad_spi_control_port_read,                      --                                                           .read
			dac_grad_spi_control_port_readdata                               => mm_interconnect_1_dac_grad_spi_control_port_readdata,                  --                                                           .readdata
			dac_grad_spi_control_port_writedata                              => mm_interconnect_1_dac_grad_spi_control_port_writedata,                 --                                                           .writedata
			dac_grad_spi_control_port_chipselect                             => mm_interconnect_1_dac_grad_spi_control_port_chipselect,                --                                                           .chipselect
			dconv_fifo_mem_in_csr_address                                    => mm_interconnect_1_dconv_fifo_mem_in_csr_address,                       --                                      dconv_fifo_mem_in_csr.address
			dconv_fifo_mem_in_csr_write                                      => mm_interconnect_1_dconv_fifo_mem_in_csr_write,                         --                                                           .write
			dconv_fifo_mem_in_csr_read                                       => mm_interconnect_1_dconv_fifo_mem_in_csr_read,                          --                                                           .read
			dconv_fifo_mem_in_csr_readdata                                   => mm_interconnect_1_dconv_fifo_mem_in_csr_readdata,                      --                                                           .readdata
			dconv_fifo_mem_in_csr_writedata                                  => mm_interconnect_1_dconv_fifo_mem_in_csr_writedata,                     --                                                           .writedata
			dconv_fifo_mem_out_address                                       => mm_interconnect_1_dconv_fifo_mem_out_address,                          --                                         dconv_fifo_mem_out.address
			dconv_fifo_mem_out_read                                          => mm_interconnect_1_dconv_fifo_mem_out_read,                             --                                                           .read
			dconv_fifo_mem_out_readdata                                      => mm_interconnect_1_dconv_fifo_mem_out_readdata,                         --                                                           .readdata
			dconv_fifo_mem_out_waitrequest                                   => mm_interconnect_1_dconv_fifo_mem_out_waitrequest,                      --                                                           .waitrequest
			dconv_fifo_mem_q_in_csr_address                                  => mm_interconnect_1_dconv_fifo_mem_q_in_csr_address,                     --                                    dconv_fifo_mem_q_in_csr.address
			dconv_fifo_mem_q_in_csr_write                                    => mm_interconnect_1_dconv_fifo_mem_q_in_csr_write,                       --                                                           .write
			dconv_fifo_mem_q_in_csr_read                                     => mm_interconnect_1_dconv_fifo_mem_q_in_csr_read,                        --                                                           .read
			dconv_fifo_mem_q_in_csr_readdata                                 => mm_interconnect_1_dconv_fifo_mem_q_in_csr_readdata,                    --                                                           .readdata
			dconv_fifo_mem_q_in_csr_writedata                                => mm_interconnect_1_dconv_fifo_mem_q_in_csr_writedata,                   --                                                           .writedata
			dconv_fifo_mem_q_out_address                                     => mm_interconnect_1_dconv_fifo_mem_q_out_address,                        --                                       dconv_fifo_mem_q_out.address
			dconv_fifo_mem_q_out_read                                        => mm_interconnect_1_dconv_fifo_mem_q_out_read,                           --                                                           .read
			dconv_fifo_mem_q_out_readdata                                    => mm_interconnect_1_dconv_fifo_mem_q_out_readdata,                       --                                                           .readdata
			dconv_fifo_mem_q_out_waitrequest                                 => mm_interconnect_1_dconv_fifo_mem_q_out_waitrequest,                    --                                                           .waitrequest
			dconv_fir_avalon_mm_slave_address                                => mm_interconnect_1_dconv_fir_avalon_mm_slave_address,                   --                                  dconv_fir_avalon_mm_slave.address
			dconv_fir_avalon_mm_slave_write                                  => mm_interconnect_1_dconv_fir_avalon_mm_slave_write,                     --                                                           .write
			dconv_fir_avalon_mm_slave_read                                   => mm_interconnect_1_dconv_fir_avalon_mm_slave_read,                      --                                                           .read
			dconv_fir_avalon_mm_slave_readdata                               => mm_interconnect_1_dconv_fir_avalon_mm_slave_readdata,                  --                                                           .readdata
			dconv_fir_avalon_mm_slave_writedata                              => mm_interconnect_1_dconv_fir_avalon_mm_slave_writedata,                 --                                                           .writedata
			dconv_fir_avalon_mm_slave_readdatavalid                          => mm_interconnect_1_dconv_fir_avalon_mm_slave_readdatavalid,             --                                                           .readdatavalid
			dconv_fir_q_avalon_mm_slave_address                              => mm_interconnect_1_dconv_fir_q_avalon_mm_slave_address,                 --                                dconv_fir_q_avalon_mm_slave.address
			dconv_fir_q_avalon_mm_slave_write                                => mm_interconnect_1_dconv_fir_q_avalon_mm_slave_write,                   --                                                           .write
			dconv_fir_q_avalon_mm_slave_read                                 => mm_interconnect_1_dconv_fir_q_avalon_mm_slave_read,                    --                                                           .read
			dconv_fir_q_avalon_mm_slave_readdata                             => mm_interconnect_1_dconv_fir_q_avalon_mm_slave_readdata,                --                                                           .readdata
			dconv_fir_q_avalon_mm_slave_writedata                            => mm_interconnect_1_dconv_fir_q_avalon_mm_slave_writedata,               --                                                           .writedata
			dconv_fir_q_avalon_mm_slave_readdatavalid                        => mm_interconnect_1_dconv_fir_q_avalon_mm_slave_readdatavalid,           --                                                           .readdatavalid
			dma_dconvi_control_port_slave_address                            => mm_interconnect_1_dma_dconvi_control_port_slave_address,               --                              dma_dconvi_control_port_slave.address
			dma_dconvi_control_port_slave_write                              => mm_interconnect_1_dma_dconvi_control_port_slave_write,                 --                                                           .write
			dma_dconvi_control_port_slave_readdata                           => mm_interconnect_1_dma_dconvi_control_port_slave_readdata,              --                                                           .readdata
			dma_dconvi_control_port_slave_writedata                          => mm_interconnect_1_dma_dconvi_control_port_slave_writedata,             --                                                           .writedata
			dma_dconvi_control_port_slave_chipselect                         => mm_interconnect_1_dma_dconvi_control_port_slave_chipselect,            --                                                           .chipselect
			dma_dconvq_control_port_slave_address                            => mm_interconnect_1_dma_dconvq_control_port_slave_address,               --                              dma_dconvq_control_port_slave.address
			dma_dconvq_control_port_slave_write                              => mm_interconnect_1_dma_dconvq_control_port_slave_write,                 --                                                           .write
			dma_dconvq_control_port_slave_readdata                           => mm_interconnect_1_dma_dconvq_control_port_slave_readdata,              --                                                           .readdata
			dma_dconvq_control_port_slave_writedata                          => mm_interconnect_1_dma_dconvq_control_port_slave_writedata,             --                                                           .writedata
			dma_dconvq_control_port_slave_chipselect                         => mm_interconnect_1_dma_dconvq_control_port_slave_chipselect,            --                                                           .chipselect
			dma_dummy_control_port_slave_address                             => mm_interconnect_1_dma_dummy_control_port_slave_address,                --                               dma_dummy_control_port_slave.address
			dma_dummy_control_port_slave_write                               => mm_interconnect_1_dma_dummy_control_port_slave_write,                  --                                                           .write
			dma_dummy_control_port_slave_readdata                            => mm_interconnect_1_dma_dummy_control_port_slave_readdata,               --                                                           .readdata
			dma_dummy_control_port_slave_writedata                           => mm_interconnect_1_dma_dummy_control_port_slave_writedata,              --                                                           .writedata
			dma_dummy_control_port_slave_chipselect                          => mm_interconnect_1_dma_dummy_control_port_slave_chipselect,             --                                                           .chipselect
			dma_fifo_control_port_slave_address                              => mm_interconnect_1_dma_fifo_control_port_slave_address,                 --                                dma_fifo_control_port_slave.address
			dma_fifo_control_port_slave_write                                => mm_interconnect_1_dma_fifo_control_port_slave_write,                   --                                                           .write
			dma_fifo_control_port_slave_readdata                             => mm_interconnect_1_dma_fifo_control_port_slave_readdata,                --                                                           .readdata
			dma_fifo_control_port_slave_writedata                            => mm_interconnect_1_dma_fifo_control_port_slave_writedata,               --                                                           .writedata
			dma_fifo_control_port_slave_chipselect                           => mm_interconnect_1_dma_fifo_control_port_slave_chipselect,              --                                                           .chipselect
			fifo_dummy_in_write                                              => mm_interconnect_1_fifo_dummy_in_write,                                 --                                              fifo_dummy_in.write
			fifo_dummy_in_writedata                                          => mm_interconnect_1_fifo_dummy_in_writedata,                             --                                                           .writedata
			fifo_dummy_in_waitrequest                                        => mm_interconnect_1_fifo_dummy_in_waitrequest,                           --                                                           .waitrequest
			fifo_dummy_in_csr_address                                        => mm_interconnect_1_fifo_dummy_in_csr_address,                           --                                          fifo_dummy_in_csr.address
			fifo_dummy_in_csr_write                                          => mm_interconnect_1_fifo_dummy_in_csr_write,                             --                                                           .write
			fifo_dummy_in_csr_read                                           => mm_interconnect_1_fifo_dummy_in_csr_read,                              --                                                           .read
			fifo_dummy_in_csr_readdata                                       => mm_interconnect_1_fifo_dummy_in_csr_readdata,                          --                                                           .readdata
			fifo_dummy_in_csr_writedata                                      => mm_interconnect_1_fifo_dummy_in_csr_writedata,                         --                                                           .writedata
			fifo_dummy_out_read                                              => mm_interconnect_1_fifo_dummy_out_read,                                 --                                             fifo_dummy_out.read
			fifo_dummy_out_readdata                                          => mm_interconnect_1_fifo_dummy_out_readdata,                             --                                                           .readdata
			fifo_dummy_out_waitrequest                                       => mm_interconnect_1_fifo_dummy_out_waitrequest,                          --                                                           .waitrequest
			fifo_dummy64_in_in_address                                       => mm_interconnect_1_fifo_dummy64_in_in_address,                          --                                         fifo_dummy64_in_in.address
			fifo_dummy64_in_in_write                                         => mm_interconnect_1_fifo_dummy64_in_in_write,                            --                                                           .write
			fifo_dummy64_in_in_writedata                                     => mm_interconnect_1_fifo_dummy64_in_in_writedata,                        --                                                           .writedata
			fifo_dummy64_in_in_waitrequest                                   => mm_interconnect_1_fifo_dummy64_in_in_waitrequest,                      --                                                           .waitrequest
			fifo_dummy64_in_in_csr_address                                   => mm_interconnect_1_fifo_dummy64_in_in_csr_address,                      --                                     fifo_dummy64_in_in_csr.address
			fifo_dummy64_in_in_csr_write                                     => mm_interconnect_1_fifo_dummy64_in_in_csr_write,                        --                                                           .write
			fifo_dummy64_in_in_csr_read                                      => mm_interconnect_1_fifo_dummy64_in_in_csr_read,                         --                                                           .read
			fifo_dummy64_in_in_csr_readdata                                  => mm_interconnect_1_fifo_dummy64_in_in_csr_readdata,                     --                                                           .readdata
			fifo_dummy64_in_in_csr_writedata                                 => mm_interconnect_1_fifo_dummy64_in_in_csr_writedata,                    --                                                           .writedata
			fifo_dummy64_out_in_csr_address                                  => mm_interconnect_1_fifo_dummy64_out_in_csr_address,                     --                                    fifo_dummy64_out_in_csr.address
			fifo_dummy64_out_in_csr_write                                    => mm_interconnect_1_fifo_dummy64_out_in_csr_write,                       --                                                           .write
			fifo_dummy64_out_in_csr_read                                     => mm_interconnect_1_fifo_dummy64_out_in_csr_read,                        --                                                           .read
			fifo_dummy64_out_in_csr_readdata                                 => mm_interconnect_1_fifo_dummy64_out_in_csr_readdata,                    --                                                           .readdata
			fifo_dummy64_out_in_csr_writedata                                => mm_interconnect_1_fifo_dummy64_out_in_csr_writedata,                   --                                                           .writedata
			fifo_dummy64_out_out_address                                     => mm_interconnect_1_fifo_dummy64_out_out_address,                        --                                       fifo_dummy64_out_out.address
			fifo_dummy64_out_out_read                                        => mm_interconnect_1_fifo_dummy64_out_out_read,                           --                                                           .read
			fifo_dummy64_out_out_readdata                                    => mm_interconnect_1_fifo_dummy64_out_out_readdata,                       --                                                           .readdata
			fifo_dummy64_out_out_waitrequest                                 => mm_interconnect_1_fifo_dummy64_out_out_waitrequest,                    --                                                           .waitrequest
			i2c_ext_csr_address                                              => mm_interconnect_1_i2c_ext_csr_address,                                 --                                                i2c_ext_csr.address
			i2c_ext_csr_write                                                => mm_interconnect_1_i2c_ext_csr_write,                                   --                                                           .write
			i2c_ext_csr_read                                                 => mm_interconnect_1_i2c_ext_csr_read,                                    --                                                           .read
			i2c_ext_csr_readdata                                             => mm_interconnect_1_i2c_ext_csr_readdata,                                --                                                           .readdata
			i2c_ext_csr_writedata                                            => mm_interconnect_1_i2c_ext_csr_writedata,                               --                                                           .writedata
			i2c_int_csr_address                                              => mm_interconnect_1_i2c_int_csr_address,                                 --                                                i2c_int_csr.address
			i2c_int_csr_write                                                => mm_interconnect_1_i2c_int_csr_write,                                   --                                                           .write
			i2c_int_csr_read                                                 => mm_interconnect_1_i2c_int_csr_read,                                    --                                                           .read
			i2c_int_csr_readdata                                             => mm_interconnect_1_i2c_int_csr_readdata,                                --                                                           .readdata
			i2c_int_csr_writedata                                            => mm_interconnect_1_i2c_int_csr_writedata,                               --                                                           .writedata
			jtag_uart_avalon_jtag_slave_address                              => mm_interconnect_1_jtag_uart_avalon_jtag_slave_address,                 --                                jtag_uart_avalon_jtag_slave.address
			jtag_uart_avalon_jtag_slave_write                                => mm_interconnect_1_jtag_uart_avalon_jtag_slave_write,                   --                                                           .write
			jtag_uart_avalon_jtag_slave_read                                 => mm_interconnect_1_jtag_uart_avalon_jtag_slave_read,                    --                                                           .read
			jtag_uart_avalon_jtag_slave_readdata                             => mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata,                --                                                           .readdata
			jtag_uart_avalon_jtag_slave_writedata                            => mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata,               --                                                           .writedata
			jtag_uart_avalon_jtag_slave_waitrequest                          => mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest,             --                                                           .waitrequest
			jtag_uart_avalon_jtag_slave_chipselect                           => mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect,              --                                                           .chipselect
			nmr_parameters_adc_val_sub_s1_address                            => mm_interconnect_1_nmr_parameters_adc_val_sub_s1_address,               --                              nmr_parameters_adc_val_sub_s1.address
			nmr_parameters_adc_val_sub_s1_write                              => mm_interconnect_1_nmr_parameters_adc_val_sub_s1_write,                 --                                                           .write
			nmr_parameters_adc_val_sub_s1_readdata                           => mm_interconnect_1_nmr_parameters_adc_val_sub_s1_readdata,              --                                                           .readdata
			nmr_parameters_adc_val_sub_s1_writedata                          => mm_interconnect_1_nmr_parameters_adc_val_sub_s1_writedata,             --                                                           .writedata
			nmr_parameters_adc_val_sub_s1_chipselect                         => mm_interconnect_1_nmr_parameters_adc_val_sub_s1_chipselect,            --                                                           .chipselect
			nmr_parameters_delay_nosig_s1_address                            => mm_interconnect_1_nmr_parameters_delay_nosig_s1_address,               --                              nmr_parameters_delay_nosig_s1.address
			nmr_parameters_delay_nosig_s1_write                              => mm_interconnect_1_nmr_parameters_delay_nosig_s1_write,                 --                                                           .write
			nmr_parameters_delay_nosig_s1_readdata                           => mm_interconnect_1_nmr_parameters_delay_nosig_s1_readdata,              --                                                           .readdata
			nmr_parameters_delay_nosig_s1_writedata                          => mm_interconnect_1_nmr_parameters_delay_nosig_s1_writedata,             --                                                           .writedata
			nmr_parameters_delay_nosig_s1_chipselect                         => mm_interconnect_1_nmr_parameters_delay_nosig_s1_chipselect,            --                                                           .chipselect
			nmr_parameters_delay_sig_s1_address                              => mm_interconnect_1_nmr_parameters_delay_sig_s1_address,                 --                                nmr_parameters_delay_sig_s1.address
			nmr_parameters_delay_sig_s1_write                                => mm_interconnect_1_nmr_parameters_delay_sig_s1_write,                   --                                                           .write
			nmr_parameters_delay_sig_s1_readdata                             => mm_interconnect_1_nmr_parameters_delay_sig_s1_readdata,                --                                                           .readdata
			nmr_parameters_delay_sig_s1_writedata                            => mm_interconnect_1_nmr_parameters_delay_sig_s1_writedata,               --                                                           .writedata
			nmr_parameters_delay_sig_s1_chipselect                           => mm_interconnect_1_nmr_parameters_delay_sig_s1_chipselect,              --                                                           .chipselect
			nmr_parameters_delay_t1_s1_address                               => mm_interconnect_1_nmr_parameters_delay_t1_s1_address,                  --                                 nmr_parameters_delay_t1_s1.address
			nmr_parameters_delay_t1_s1_write                                 => mm_interconnect_1_nmr_parameters_delay_t1_s1_write,                    --                                                           .write
			nmr_parameters_delay_t1_s1_readdata                              => mm_interconnect_1_nmr_parameters_delay_t1_s1_readdata,                 --                                                           .readdata
			nmr_parameters_delay_t1_s1_writedata                             => mm_interconnect_1_nmr_parameters_delay_t1_s1_writedata,                --                                                           .writedata
			nmr_parameters_delay_t1_s1_chipselect                            => mm_interconnect_1_nmr_parameters_delay_t1_s1_chipselect,               --                                                           .chipselect
			nmr_parameters_echoes_per_scan_s1_address                        => mm_interconnect_1_nmr_parameters_echoes_per_scan_s1_address,           --                          nmr_parameters_echoes_per_scan_s1.address
			nmr_parameters_echoes_per_scan_s1_write                          => mm_interconnect_1_nmr_parameters_echoes_per_scan_s1_write,             --                                                           .write
			nmr_parameters_echoes_per_scan_s1_readdata                       => mm_interconnect_1_nmr_parameters_echoes_per_scan_s1_readdata,          --                                                           .readdata
			nmr_parameters_echoes_per_scan_s1_writedata                      => mm_interconnect_1_nmr_parameters_echoes_per_scan_s1_writedata,         --                                                           .writedata
			nmr_parameters_echoes_per_scan_s1_chipselect                     => mm_interconnect_1_nmr_parameters_echoes_per_scan_s1_chipselect,        --                                                           .chipselect
			nmr_parameters_init_delay_s1_address                             => mm_interconnect_1_nmr_parameters_init_delay_s1_address,                --                               nmr_parameters_init_delay_s1.address
			nmr_parameters_init_delay_s1_write                               => mm_interconnect_1_nmr_parameters_init_delay_s1_write,                  --                                                           .write
			nmr_parameters_init_delay_s1_readdata                            => mm_interconnect_1_nmr_parameters_init_delay_s1_readdata,               --                                                           .readdata
			nmr_parameters_init_delay_s1_writedata                           => mm_interconnect_1_nmr_parameters_init_delay_s1_writedata,              --                                                           .writedata
			nmr_parameters_init_delay_s1_chipselect                          => mm_interconnect_1_nmr_parameters_init_delay_s1_chipselect,             --                                                           .chipselect
			nmr_parameters_pulse_180deg_s1_address                           => mm_interconnect_1_nmr_parameters_pulse_180deg_s1_address,              --                             nmr_parameters_pulse_180deg_s1.address
			nmr_parameters_pulse_180deg_s1_write                             => mm_interconnect_1_nmr_parameters_pulse_180deg_s1_write,                --                                                           .write
			nmr_parameters_pulse_180deg_s1_readdata                          => mm_interconnect_1_nmr_parameters_pulse_180deg_s1_readdata,             --                                                           .readdata
			nmr_parameters_pulse_180deg_s1_writedata                         => mm_interconnect_1_nmr_parameters_pulse_180deg_s1_writedata,            --                                                           .writedata
			nmr_parameters_pulse_180deg_s1_chipselect                        => mm_interconnect_1_nmr_parameters_pulse_180deg_s1_chipselect,           --                                                           .chipselect
			nmr_parameters_pulse_90deg_s1_address                            => mm_interconnect_1_nmr_parameters_pulse_90deg_s1_address,               --                              nmr_parameters_pulse_90deg_s1.address
			nmr_parameters_pulse_90deg_s1_write                              => mm_interconnect_1_nmr_parameters_pulse_90deg_s1_write,                 --                                                           .write
			nmr_parameters_pulse_90deg_s1_readdata                           => mm_interconnect_1_nmr_parameters_pulse_90deg_s1_readdata,              --                                                           .readdata
			nmr_parameters_pulse_90deg_s1_writedata                          => mm_interconnect_1_nmr_parameters_pulse_90deg_s1_writedata,             --                                                           .writedata
			nmr_parameters_pulse_90deg_s1_chipselect                         => mm_interconnect_1_nmr_parameters_pulse_90deg_s1_chipselect,            --                                                           .chipselect
			nmr_parameters_pulse_t1_s1_address                               => mm_interconnect_1_nmr_parameters_pulse_t1_s1_address,                  --                                 nmr_parameters_pulse_t1_s1.address
			nmr_parameters_pulse_t1_s1_write                                 => mm_interconnect_1_nmr_parameters_pulse_t1_s1_write,                    --                                                           .write
			nmr_parameters_pulse_t1_s1_readdata                              => mm_interconnect_1_nmr_parameters_pulse_t1_s1_readdata,                 --                                                           .readdata
			nmr_parameters_pulse_t1_s1_writedata                             => mm_interconnect_1_nmr_parameters_pulse_t1_s1_writedata,                --                                                           .writedata
			nmr_parameters_pulse_t1_s1_chipselect                            => mm_interconnect_1_nmr_parameters_pulse_t1_s1_chipselect,               --                                                           .chipselect
			nmr_parameters_rx_delay_s1_address                               => mm_interconnect_1_nmr_parameters_rx_delay_s1_address,                  --                                 nmr_parameters_rx_delay_s1.address
			nmr_parameters_rx_delay_s1_write                                 => mm_interconnect_1_nmr_parameters_rx_delay_s1_write,                    --                                                           .write
			nmr_parameters_rx_delay_s1_readdata                              => mm_interconnect_1_nmr_parameters_rx_delay_s1_readdata,                 --                                                           .readdata
			nmr_parameters_rx_delay_s1_writedata                             => mm_interconnect_1_nmr_parameters_rx_delay_s1_writedata,                --                                                           .writedata
			nmr_parameters_rx_delay_s1_chipselect                            => mm_interconnect_1_nmr_parameters_rx_delay_s1_chipselect,               --                                                           .chipselect
			nmr_parameters_samples_per_echo_s1_address                       => mm_interconnect_1_nmr_parameters_samples_per_echo_s1_address,          --                         nmr_parameters_samples_per_echo_s1.address
			nmr_parameters_samples_per_echo_s1_write                         => mm_interconnect_1_nmr_parameters_samples_per_echo_s1_write,            --                                                           .write
			nmr_parameters_samples_per_echo_s1_readdata                      => mm_interconnect_1_nmr_parameters_samples_per_echo_s1_readdata,         --                                                           .readdata
			nmr_parameters_samples_per_echo_s1_writedata                     => mm_interconnect_1_nmr_parameters_samples_per_echo_s1_writedata,        --                                                           .writedata
			nmr_parameters_samples_per_echo_s1_chipselect                    => mm_interconnect_1_nmr_parameters_samples_per_echo_s1_chipselect,       --                                                           .chipselect
			nmr_sys_pll_reconfig_mgmt_avalon_slave_address                   => mm_interconnect_1_nmr_sys_pll_reconfig_mgmt_avalon_slave_address,      --                     nmr_sys_pll_reconfig_mgmt_avalon_slave.address
			nmr_sys_pll_reconfig_mgmt_avalon_slave_write                     => mm_interconnect_1_nmr_sys_pll_reconfig_mgmt_avalon_slave_write,        --                                                           .write
			nmr_sys_pll_reconfig_mgmt_avalon_slave_read                      => mm_interconnect_1_nmr_sys_pll_reconfig_mgmt_avalon_slave_read,         --                                                           .read
			nmr_sys_pll_reconfig_mgmt_avalon_slave_readdata                  => mm_interconnect_1_nmr_sys_pll_reconfig_mgmt_avalon_slave_readdata,     --                                                           .readdata
			nmr_sys_pll_reconfig_mgmt_avalon_slave_writedata                 => mm_interconnect_1_nmr_sys_pll_reconfig_mgmt_avalon_slave_writedata,    --                                                           .writedata
			nmr_sys_pll_reconfig_mgmt_avalon_slave_waitrequest               => mm_interconnect_1_nmr_sys_pll_reconfig_mgmt_avalon_slave_waitrequest,  --                                                           .waitrequest
			sdram_s1_address                                                 => mm_interconnect_1_sdram_s1_address,                                    --                                                   sdram_s1.address
			sdram_s1_write                                                   => mm_interconnect_1_sdram_s1_write,                                      --                                                           .write
			sdram_s1_read                                                    => mm_interconnect_1_sdram_s1_read,                                       --                                                           .read
			sdram_s1_readdata                                                => mm_interconnect_1_sdram_s1_readdata,                                   --                                                           .readdata
			sdram_s1_writedata                                               => mm_interconnect_1_sdram_s1_writedata,                                  --                                                           .writedata
			sdram_s1_byteenable                                              => mm_interconnect_1_sdram_s1_byteenable,                                 --                                                           .byteenable
			sdram_s1_readdatavalid                                           => mm_interconnect_1_sdram_s1_readdatavalid,                              --                                                           .readdatavalid
			sdram_s1_waitrequest                                             => mm_interconnect_1_sdram_s1_waitrequest,                                --                                                           .waitrequest
			sdram_s1_chipselect                                              => mm_interconnect_1_sdram_s1_chipselect,                                 --                                                           .chipselect
			spi_afe_relays_spi_control_port_address                          => mm_interconnect_1_spi_afe_relays_spi_control_port_address,             --                            spi_afe_relays_spi_control_port.address
			spi_afe_relays_spi_control_port_write                            => mm_interconnect_1_spi_afe_relays_spi_control_port_write,               --                                                           .write
			spi_afe_relays_spi_control_port_read                             => mm_interconnect_1_spi_afe_relays_spi_control_port_read,                --                                                           .read
			spi_afe_relays_spi_control_port_readdata                         => mm_interconnect_1_spi_afe_relays_spi_control_port_readdata,            --                                                           .readdata
			spi_afe_relays_spi_control_port_writedata                        => mm_interconnect_1_spi_afe_relays_spi_control_port_writedata,           --                                                           .writedata
			spi_afe_relays_spi_control_port_chipselect                       => mm_interconnect_1_spi_afe_relays_spi_control_port_chipselect,          --                                                           .chipselect
			spi_mtch_ntwrk_spi_control_port_address                          => mm_interconnect_1_spi_mtch_ntwrk_spi_control_port_address,             --                            spi_mtch_ntwrk_spi_control_port.address
			spi_mtch_ntwrk_spi_control_port_write                            => mm_interconnect_1_spi_mtch_ntwrk_spi_control_port_write,               --                                                           .write
			spi_mtch_ntwrk_spi_control_port_read                             => mm_interconnect_1_spi_mtch_ntwrk_spi_control_port_read,                --                                                           .read
			spi_mtch_ntwrk_spi_control_port_readdata                         => mm_interconnect_1_spi_mtch_ntwrk_spi_control_port_readdata,            --                                                           .readdata
			spi_mtch_ntwrk_spi_control_port_writedata                        => mm_interconnect_1_spi_mtch_ntwrk_spi_control_port_writedata,           --                                                           .writedata
			spi_mtch_ntwrk_spi_control_port_chipselect                       => mm_interconnect_1_spi_mtch_ntwrk_spi_control_port_chipselect,          --                                                           .chipselect
			switches_s1_address                                              => mm_interconnect_1_switches_s1_address,                                 --                                                switches_s1.address
			switches_s1_readdata                                             => mm_interconnect_1_switches_s1_readdata,                                --                                                           .readdata
			sysid_qsys_control_slave_address                                 => mm_interconnect_1_sysid_qsys_control_slave_address,                    --                                   sysid_qsys_control_slave.address
			sysid_qsys_control_slave_readdata                                => mm_interconnect_1_sysid_qsys_control_slave_readdata                    --                                                           .readdata
		);

	irq_mapper : component soc_system_v5_irq_mapper
		port map (
			clk           => open,                     --       clk.clk
			reset         => open,                     -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq, -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq, -- receiver1.irq
			sender_irq    => hps_0_f2h_irq0_irq        --    sender.irq
		);

	irq_mapper_001 : component soc_system_v5_irq_mapper_001
		port map (
			clk           => open,                         --       clk.clk
			reset         => open,                         -- clk_reset.reset
			receiver0_irq => irq_mapper_001_receiver0_irq, -- receiver0.irq
			receiver1_irq => irq_mapper_001_receiver1_irq, -- receiver1.irq
			receiver2_irq => irq_mapper_001_receiver2_irq, -- receiver2.irq
			receiver3_irq => irq_mapper_001_receiver3_irq, -- receiver3.irq
			receiver4_irq => irq_mapper_001_receiver4_irq, -- receiver4.irq
			receiver5_irq => irq_mapper_001_receiver5_irq, -- receiver5.irq
			receiver6_irq => irq_mapper_001_receiver6_irq, -- receiver6.irq
			receiver7_irq => irq_mapper_001_receiver7_irq, -- receiver7.irq
			sender_irq    => hps_0_f2h_irq1_irq            --    sender.irq
		);

	avalon_st_adapter : component soc_system_v5_avalon_st_adapter
		generic map (
			inBitsPerSymbol => 16,
			inUsePackets    => 0,
			inDataWidth     => 16,
			inChannelWidth  => 0,
			inErrorWidth    => 0,
			inUseEmptyPort  => 0,
			inUseValid      => 1,
			inUseReady      => 1,
			inReadyLatency  => 0,
			outDataWidth    => 32,
			outChannelWidth => 0,
			outErrorWidth   => 0,
			outUseEmptyPort => 0,
			outUseValid     => 1,
			outUseReady     => 1,
			outReadyLatency => 1
		)
		port map (
			in_clk_0_clk   => clk_clk,                            -- in_clk_0.clk
			in_rst_0_reset => rst_controller_001_reset_out_reset, -- in_rst_0.reset
			in_0_data      => adc_fifo_dc_out_data,               --     in_0.data
			in_0_valid     => adc_fifo_dc_out_valid,              --         .valid
			in_0_ready     => adc_fifo_dc_out_ready,              --         .ready
			out_0_data     => avalon_st_adapter_out_0_data,       --    out_0.data
			out_0_valid    => avalon_st_adapter_out_0_valid,      --         .valid
			out_0_ready    => avalon_st_adapter_out_0_ready       --         .ready
		);

	avalon_st_adapter_001 : component soc_system_v5_avalon_st_adapter_001
		generic map (
			inBitsPerSymbol => 32,
			inUsePackets    => 0,
			inDataWidth     => 32,
			inChannelWidth  => 0,
			inErrorWidth    => 0,
			inUseEmptyPort  => 0,
			inUseValid      => 1,
			inUseReady      => 1,
			inReadyLatency  => 0,
			outDataWidth    => 32,
			outChannelWidth => 0,
			outErrorWidth   => 0,
			outUseEmptyPort => 0,
			outUseValid     => 1,
			outUseReady     => 1,
			outReadyLatency => 1
		)
		port map (
			in_clk_0_clk   => clk_clk,                            -- in_clk_0.clk
			in_rst_0_reset => rst_controller_001_reset_out_reset, -- in_rst_0.reset
			in_0_data      => dconv_fifo_dc_out_data,             --     in_0.data
			in_0_valid     => dconv_fifo_dc_out_valid,            --         .valid
			in_0_ready     => dconv_fifo_dc_out_ready,            --         .ready
			out_0_data     => avalon_st_adapter_001_out_0_data,   --    out_0.data
			out_0_valid    => avalon_st_adapter_001_out_0_valid,  --         .valid
			out_0_ready    => avalon_st_adapter_001_out_0_ready   --         .ready
		);

	avalon_st_adapter_002 : component soc_system_v5_avalon_st_adapter_001
		generic map (
			inBitsPerSymbol => 32,
			inUsePackets    => 0,
			inDataWidth     => 32,
			inChannelWidth  => 0,
			inErrorWidth    => 0,
			inUseEmptyPort  => 0,
			inUseValid      => 1,
			inUseReady      => 1,
			inReadyLatency  => 0,
			outDataWidth    => 32,
			outChannelWidth => 0,
			outErrorWidth   => 0,
			outUseEmptyPort => 0,
			outUseValid     => 1,
			outUseReady     => 1,
			outReadyLatency => 1
		)
		port map (
			in_clk_0_clk   => clk_clk,                            -- in_clk_0.clk
			in_rst_0_reset => rst_controller_001_reset_out_reset, -- in_rst_0.reset
			in_0_data      => dconv_fifo_dc_q_out_data,           --     in_0.data
			in_0_valid     => dconv_fifo_dc_q_out_valid,          --         .valid
			in_0_ready     => dconv_fifo_dc_q_out_ready,          --         .ready
			out_0_data     => avalon_st_adapter_002_out_0_data,   --    out_0.data
			out_0_valid    => avalon_st_adapter_002_out_0_valid,  --         .valid
			out_0_ready    => avalon_st_adapter_002_out_0_ready   --         .ready
		);

	rst_controller : component soc_system_v5_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,        -- reset_in0.reset
			reset_in1      => fifo_rst_reset,                 -- reset_in1.reset
			clk            => fifo_clk_bridge_in_clk,         --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	rst_controller_001 : component soc_system_v5_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => fifo_rst_reset,                     -- reset_in1.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_002 : component soc_system_v5_rst_controller_002
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => gp_pll_outclk0_clk,                 --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_003 : component soc_system_v5_rst_controller_002
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_003_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_004 : component soc_system_v5_rst_controller_002
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => hps_0_h2f_reset_reset_n_ports_inv,  -- reset_in0.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_004_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	fifo_rst_reset_ports_inv <= not fifo_rst_reset;

	hps_0_h2f_reset_reset_n_ports_inv <= not hps_0_h2f_reset_reset;

	reset_reset_n_ports_inv <= not reset_reset_n;

	dma_fifo_write_master_write_ports_inv <= not dma_fifo_write_master_write;

	dma_dconvi_write_master_write_ports_inv <= not dma_dconvi_write_master_write;

	dma_dconvq_write_master_write_ports_inv <= not dma_dconvq_write_master_write;

	dma_dummy_write_master_write_ports_inv <= not dma_dummy_write_master_write;

	dma_fifo_read_master_read_ports_inv <= not dma_fifo_read_master_read;

	dma_dconvq_read_master_read_ports_inv <= not dma_dconvq_read_master_read;

	dma_dconvi_read_master_read_ports_inv <= not dma_dconvi_read_master_read;

	dma_dummy_read_master_read_ports_inv <= not dma_dummy_read_master_read;

	mm_interconnect_1_sdram_s1_read_ports_inv <= not mm_interconnect_1_sdram_s1_read;

	mm_interconnect_1_sdram_s1_byteenable_ports_inv <= not mm_interconnect_1_sdram_s1_byteenable;

	mm_interconnect_1_sdram_s1_write_ports_inv <= not mm_interconnect_1_sdram_s1_write;

	mm_interconnect_1_nmr_parameters_adc_val_sub_s1_write_ports_inv <= not mm_interconnect_1_nmr_parameters_adc_val_sub_s1_write;

	mm_interconnect_1_jtag_uart_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_1_jtag_uart_avalon_jtag_slave_read;

	mm_interconnect_1_jtag_uart_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_1_jtag_uart_avalon_jtag_slave_write;

	mm_interconnect_1_nmr_parameters_delay_nosig_s1_write_ports_inv <= not mm_interconnect_1_nmr_parameters_delay_nosig_s1_write;

	mm_interconnect_1_nmr_parameters_delay_sig_s1_write_ports_inv <= not mm_interconnect_1_nmr_parameters_delay_sig_s1_write;

	mm_interconnect_1_nmr_parameters_delay_t1_s1_write_ports_inv <= not mm_interconnect_1_nmr_parameters_delay_t1_s1_write;

	mm_interconnect_1_nmr_parameters_echoes_per_scan_s1_write_ports_inv <= not mm_interconnect_1_nmr_parameters_echoes_per_scan_s1_write;

	mm_interconnect_1_nmr_parameters_init_delay_s1_write_ports_inv <= not mm_interconnect_1_nmr_parameters_init_delay_s1_write;

	mm_interconnect_1_nmr_parameters_pulse_180deg_s1_write_ports_inv <= not mm_interconnect_1_nmr_parameters_pulse_180deg_s1_write;

	mm_interconnect_1_nmr_parameters_pulse_90deg_s1_write_ports_inv <= not mm_interconnect_1_nmr_parameters_pulse_90deg_s1_write;

	mm_interconnect_1_nmr_parameters_pulse_t1_s1_write_ports_inv <= not mm_interconnect_1_nmr_parameters_pulse_t1_s1_write;

	mm_interconnect_1_nmr_parameters_rx_delay_s1_write_ports_inv <= not mm_interconnect_1_nmr_parameters_rx_delay_s1_write;

	mm_interconnect_1_ctrl_out_s1_write_ports_inv <= not mm_interconnect_1_ctrl_out_s1_write;

	mm_interconnect_1_aux_cnt_out_s1_write_ports_inv <= not mm_interconnect_1_aux_cnt_out_s1_write;

	mm_interconnect_1_nmr_parameters_samples_per_echo_s1_write_ports_inv <= not mm_interconnect_1_nmr_parameters_samples_per_echo_s1_write;

	mm_interconnect_1_dac_grad_spi_control_port_read_ports_inv <= not mm_interconnect_1_dac_grad_spi_control_port_read;

	mm_interconnect_1_dac_grad_spi_control_port_write_ports_inv <= not mm_interconnect_1_dac_grad_spi_control_port_write;

	mm_interconnect_1_spi_mtch_ntwrk_spi_control_port_read_ports_inv <= not mm_interconnect_1_spi_mtch_ntwrk_spi_control_port_read;

	mm_interconnect_1_spi_mtch_ntwrk_spi_control_port_write_ports_inv <= not mm_interconnect_1_spi_mtch_ntwrk_spi_control_port_write;

	mm_interconnect_1_spi_afe_relays_spi_control_port_read_ports_inv <= not mm_interconnect_1_spi_afe_relays_spi_control_port_read;

	mm_interconnect_1_spi_afe_relays_spi_control_port_write_ports_inv <= not mm_interconnect_1_spi_afe_relays_spi_control_port_write;

	mm_interconnect_1_dma_fifo_control_port_slave_write_ports_inv <= not mm_interconnect_1_dma_fifo_control_port_slave_write;

	mm_interconnect_1_dma_dconvi_control_port_slave_write_ports_inv <= not mm_interconnect_1_dma_dconvi_control_port_slave_write;

	mm_interconnect_1_dma_dconvq_control_port_slave_write_ports_inv <= not mm_interconnect_1_dma_dconvq_control_port_slave_write;

	mm_interconnect_1_dma_dummy_control_port_slave_write_ports_inv <= not mm_interconnect_1_dma_dummy_control_port_slave_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

	rst_controller_003_reset_out_reset_ports_inv <= not rst_controller_003_reset_out_reset;

	hps_0_h2f_reset_reset_n <= hps_0_h2f_reset_reset;

end architecture rtl; -- of soc_system_v5
