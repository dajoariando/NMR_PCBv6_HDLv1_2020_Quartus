// system_parameters_0.v

// Generated using ACDS version 17.1 590

`timescale 1 ps / 1 ps
module system_parameters_0 (
		input  wire        clk_clk,                                     //                                  clk.clk
		output wire [31:0] delay_nosig_external_connection_export,      //      delay_nosig_external_connection.export
		input  wire [1:0]  delay_nosig_s1_address,                      //                       delay_nosig_s1.address
		input  wire        delay_nosig_s1_write_n,                      //                                     .write_n
		input  wire [31:0] delay_nosig_s1_writedata,                    //                                     .writedata
		input  wire        delay_nosig_s1_chipselect,                   //                                     .chipselect
		output wire [31:0] delay_nosig_s1_readdata,                     //                                     .readdata
		output wire [31:0] delay_sig_external_connection_export,        //        delay_sig_external_connection.export
		input  wire [1:0]  delay_sig_s1_address,                        //                         delay_sig_s1.address
		input  wire        delay_sig_s1_write_n,                        //                                     .write_n
		input  wire [31:0] delay_sig_s1_writedata,                      //                                     .writedata
		input  wire        delay_sig_s1_chipselect,                     //                                     .chipselect
		output wire [31:0] delay_sig_s1_readdata,                       //                                     .readdata
		output wire [31:0] delay_t1_external_connection_export,         //         delay_t1_external_connection.export
		input  wire [1:0]  delay_t1_s1_address,                         //                          delay_t1_s1.address
		input  wire        delay_t1_s1_write_n,                         //                                     .write_n
		input  wire [31:0] delay_t1_s1_writedata,                       //                                     .writedata
		input  wire        delay_t1_s1_chipselect,                      //                                     .chipselect
		output wire [31:0] delay_t1_s1_readdata,                        //                                     .readdata
		output wire [31:0] echoes_per_scan_external_connection_export,  //  echoes_per_scan_external_connection.export
		input  wire [1:0]  echoes_per_scan_s1_address,                  //                   echoes_per_scan_s1.address
		input  wire        echoes_per_scan_s1_write_n,                  //                                     .write_n
		input  wire [31:0] echoes_per_scan_s1_writedata,                //                                     .writedata
		input  wire        echoes_per_scan_s1_chipselect,               //                                     .chipselect
		output wire [31:0] echoes_per_scan_s1_readdata,                 //                                     .readdata
		output wire [31:0] init_delay_external_connection_export,       //       init_delay_external_connection.export
		input  wire [1:0]  init_delay_s1_address,                       //                        init_delay_s1.address
		input  wire        init_delay_s1_write_n,                       //                                     .write_n
		input  wire [31:0] init_delay_s1_writedata,                     //                                     .writedata
		input  wire        init_delay_s1_chipselect,                    //                                     .chipselect
		output wire [31:0] init_delay_s1_readdata,                      //                                     .readdata
		output wire [31:0] pulse_180deg_external_connection_export,     //     pulse_180deg_external_connection.export
		input  wire [1:0]  pulse_180deg_s1_address,                     //                      pulse_180deg_s1.address
		input  wire        pulse_180deg_s1_write_n,                     //                                     .write_n
		input  wire [31:0] pulse_180deg_s1_writedata,                   //                                     .writedata
		input  wire        pulse_180deg_s1_chipselect,                  //                                     .chipselect
		output wire [31:0] pulse_180deg_s1_readdata,                    //                                     .readdata
		output wire [31:0] pulse_90deg_external_connection_export,      //      pulse_90deg_external_connection.export
		input  wire [1:0]  pulse_90deg_s1_address,                      //                       pulse_90deg_s1.address
		input  wire        pulse_90deg_s1_write_n,                      //                                     .write_n
		input  wire [31:0] pulse_90deg_s1_writedata,                    //                                     .writedata
		input  wire        pulse_90deg_s1_chipselect,                   //                                     .chipselect
		output wire [31:0] pulse_90deg_s1_readdata,                     //                                     .readdata
		output wire [31:0] pulse_t1_external_connection_export,         //         pulse_t1_external_connection.export
		input  wire [1:0]  pulse_t1_s1_address,                         //                          pulse_t1_s1.address
		input  wire        pulse_t1_s1_write_n,                         //                                     .write_n
		input  wire [31:0] pulse_t1_s1_writedata,                       //                                     .writedata
		input  wire        pulse_t1_s1_chipselect,                      //                                     .chipselect
		output wire [31:0] pulse_t1_s1_readdata,                        //                                     .readdata
		input  wire        reset_reset_n,                               //                                reset.reset_n
		output wire [31:0] samples_per_echo_external_connection_export, // samples_per_echo_external_connection.export
		input  wire [1:0]  samples_per_echo_s1_address,                 //                  samples_per_echo_s1.address
		input  wire        samples_per_echo_s1_write_n,                 //                                     .write_n
		input  wire [31:0] samples_per_echo_s1_writedata,               //                                     .writedata
		input  wire        samples_per_echo_s1_chipselect,              //                                     .chipselect
		output wire [31:0] samples_per_echo_s1_readdata                 //                                     .readdata
	);

	wire    rst_controller_reset_out_reset; // rst_controller:reset_out -> [delay_nosig:reset_n, delay_sig:reset_n, delay_t1:reset_n, echoes_per_scan:reset_n, init_delay:reset_n, pulse_180deg:reset_n, pulse_90deg:reset_n, pulse_t1:reset_n, samples_per_echo:reset_n]

	system_parameters_0_delay_nosig delay_nosig (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (delay_nosig_s1_address),                 //                  s1.address
		.write_n    (delay_nosig_s1_write_n),                 //                    .write_n
		.writedata  (delay_nosig_s1_writedata),               //                    .writedata
		.chipselect (delay_nosig_s1_chipselect),              //                    .chipselect
		.readdata   (delay_nosig_s1_readdata),                //                    .readdata
		.out_port   (delay_nosig_external_connection_export)  // external_connection.export
	);

	system_parameters_0_delay_nosig delay_sig (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (delay_sig_s1_address),                 //                  s1.address
		.write_n    (delay_sig_s1_write_n),                 //                    .write_n
		.writedata  (delay_sig_s1_writedata),               //                    .writedata
		.chipselect (delay_sig_s1_chipselect),              //                    .chipselect
		.readdata   (delay_sig_s1_readdata),                //                    .readdata
		.out_port   (delay_sig_external_connection_export)  // external_connection.export
	);

	system_parameters_0_delay_t1 delay_t1 (
		.clk        (clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (delay_t1_s1_address),                 //                  s1.address
		.write_n    (delay_t1_s1_write_n),                 //                    .write_n
		.writedata  (delay_t1_s1_writedata),               //                    .writedata
		.chipselect (delay_t1_s1_chipselect),              //                    .chipselect
		.readdata   (delay_t1_s1_readdata),                //                    .readdata
		.out_port   (delay_t1_external_connection_export)  // external_connection.export
	);

	system_parameters_0_delay_t1 echoes_per_scan (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (echoes_per_scan_s1_address),                 //                  s1.address
		.write_n    (echoes_per_scan_s1_write_n),                 //                    .write_n
		.writedata  (echoes_per_scan_s1_writedata),               //                    .writedata
		.chipselect (echoes_per_scan_s1_chipselect),              //                    .chipselect
		.readdata   (echoes_per_scan_s1_readdata),                //                    .readdata
		.out_port   (echoes_per_scan_external_connection_export)  // external_connection.export
	);

	system_parameters_0_delay_t1 init_delay (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (init_delay_s1_address),                 //                  s1.address
		.write_n    (init_delay_s1_write_n),                 //                    .write_n
		.writedata  (init_delay_s1_writedata),               //                    .writedata
		.chipselect (init_delay_s1_chipselect),              //                    .chipselect
		.readdata   (init_delay_s1_readdata),                //                    .readdata
		.out_port   (init_delay_external_connection_export)  // external_connection.export
	);

	system_parameters_0_delay_nosig pulse_180deg (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (pulse_180deg_s1_address),                 //                  s1.address
		.write_n    (pulse_180deg_s1_write_n),                 //                    .write_n
		.writedata  (pulse_180deg_s1_writedata),               //                    .writedata
		.chipselect (pulse_180deg_s1_chipselect),              //                    .chipselect
		.readdata   (pulse_180deg_s1_readdata),                //                    .readdata
		.out_port   (pulse_180deg_external_connection_export)  // external_connection.export
	);

	system_parameters_0_delay_nosig pulse_90deg (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (pulse_90deg_s1_address),                 //                  s1.address
		.write_n    (pulse_90deg_s1_write_n),                 //                    .write_n
		.writedata  (pulse_90deg_s1_writedata),               //                    .writedata
		.chipselect (pulse_90deg_s1_chipselect),              //                    .chipselect
		.readdata   (pulse_90deg_s1_readdata),                //                    .readdata
		.out_port   (pulse_90deg_external_connection_export)  // external_connection.export
	);

	system_parameters_0_delay_t1 pulse_t1 (
		.clk        (clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (pulse_t1_s1_address),                 //                  s1.address
		.write_n    (pulse_t1_s1_write_n),                 //                    .write_n
		.writedata  (pulse_t1_s1_writedata),               //                    .writedata
		.chipselect (pulse_t1_s1_chipselect),              //                    .chipselect
		.readdata   (pulse_t1_s1_readdata),                //                    .readdata
		.out_port   (pulse_t1_external_connection_export)  // external_connection.export
	);

	system_parameters_0_samples_per_echo samples_per_echo (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (samples_per_echo_s1_address),                 //                  s1.address
		.write_n    (samples_per_echo_s1_write_n),                 //                    .write_n
		.writedata  (samples_per_echo_s1_writedata),               //                    .writedata
		.chipselect (samples_per_echo_s1_chipselect),              //                    .chipselect
		.readdata   (samples_per_echo_s1_readdata),                //                    .readdata
		.out_port   (samples_per_echo_external_connection_export)  // external_connection.export
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
