// soc_system_v5_nmr_parameters.v

// Generated using ACDS version 17.1 590

`timescale 1 ps / 1 ps
module soc_system_v5_nmr_parameters (
		input  wire        adc_val_sub_clk_clk,                         //                      adc_val_sub_clk.clk
		output wire [31:0] adc_val_sub_external_connection_export,      //      adc_val_sub_external_connection.export
		input  wire        adc_val_sub_reset_reset_n,                   //                    adc_val_sub_reset.reset_n
		input  wire [1:0]  adc_val_sub_s1_address,                      //                       adc_val_sub_s1.address
		input  wire        adc_val_sub_s1_write_n,                      //                                     .write_n
		input  wire [31:0] adc_val_sub_s1_writedata,                    //                                     .writedata
		input  wire        adc_val_sub_s1_chipselect,                   //                                     .chipselect
		output wire [31:0] adc_val_sub_s1_readdata,                     //                                     .readdata
		input  wire        delay_nosig_clk_clk,                         //                      delay_nosig_clk.clk
		output wire [31:0] delay_nosig_external_connection_export,      //      delay_nosig_external_connection.export
		input  wire        delay_nosig_reset_reset_n,                   //                    delay_nosig_reset.reset_n
		input  wire [1:0]  delay_nosig_s1_address,                      //                       delay_nosig_s1.address
		input  wire        delay_nosig_s1_write_n,                      //                                     .write_n
		input  wire [31:0] delay_nosig_s1_writedata,                    //                                     .writedata
		input  wire        delay_nosig_s1_chipselect,                   //                                     .chipselect
		output wire [31:0] delay_nosig_s1_readdata,                     //                                     .readdata
		input  wire        delay_sig_clk_clk,                           //                        delay_sig_clk.clk
		output wire [31:0] delay_sig_external_connection_export,        //        delay_sig_external_connection.export
		input  wire        delay_sig_reset_reset_n,                     //                      delay_sig_reset.reset_n
		input  wire [1:0]  delay_sig_s1_address,                        //                         delay_sig_s1.address
		input  wire        delay_sig_s1_write_n,                        //                                     .write_n
		input  wire [31:0] delay_sig_s1_writedata,                      //                                     .writedata
		input  wire        delay_sig_s1_chipselect,                     //                                     .chipselect
		output wire [31:0] delay_sig_s1_readdata,                       //                                     .readdata
		input  wire        delay_t1_clk_clk,                            //                         delay_t1_clk.clk
		output wire [31:0] delay_t1_external_connection_export,         //         delay_t1_external_connection.export
		input  wire        delay_t1_reset_reset_n,                      //                       delay_t1_reset.reset_n
		input  wire [1:0]  delay_t1_s1_address,                         //                          delay_t1_s1.address
		input  wire        delay_t1_s1_write_n,                         //                                     .write_n
		input  wire [31:0] delay_t1_s1_writedata,                       //                                     .writedata
		input  wire        delay_t1_s1_chipselect,                      //                                     .chipselect
		output wire [31:0] delay_t1_s1_readdata,                        //                                     .readdata
		input  wire        echoes_per_scan_clk_clk,                     //                  echoes_per_scan_clk.clk
		output wire [31:0] echoes_per_scan_external_connection_export,  //  echoes_per_scan_external_connection.export
		input  wire        echoes_per_scan_reset_reset_n,               //                echoes_per_scan_reset.reset_n
		input  wire [1:0]  echoes_per_scan_s1_address,                  //                   echoes_per_scan_s1.address
		input  wire        echoes_per_scan_s1_write_n,                  //                                     .write_n
		input  wire [31:0] echoes_per_scan_s1_writedata,                //                                     .writedata
		input  wire        echoes_per_scan_s1_chipselect,               //                                     .chipselect
		output wire [31:0] echoes_per_scan_s1_readdata,                 //                                     .readdata
		input  wire        init_delay_clk_clk,                          //                       init_delay_clk.clk
		output wire [31:0] init_delay_external_connection_export,       //       init_delay_external_connection.export
		input  wire        init_delay_reset_reset_n,                    //                     init_delay_reset.reset_n
		input  wire [1:0]  init_delay_s1_address,                       //                        init_delay_s1.address
		input  wire        init_delay_s1_write_n,                       //                                     .write_n
		input  wire [31:0] init_delay_s1_writedata,                     //                                     .writedata
		input  wire        init_delay_s1_chipselect,                    //                                     .chipselect
		output wire [31:0] init_delay_s1_readdata,                      //                                     .readdata
		input  wire        pulse_180deg_clk_clk,                        //                     pulse_180deg_clk.clk
		output wire [31:0] pulse_180deg_external_connection_export,     //     pulse_180deg_external_connection.export
		input  wire        pulse_180deg_reset_reset_n,                  //                   pulse_180deg_reset.reset_n
		input  wire [1:0]  pulse_180deg_s1_address,                     //                      pulse_180deg_s1.address
		input  wire        pulse_180deg_s1_write_n,                     //                                     .write_n
		input  wire [31:0] pulse_180deg_s1_writedata,                   //                                     .writedata
		input  wire        pulse_180deg_s1_chipselect,                  //                                     .chipselect
		output wire [31:0] pulse_180deg_s1_readdata,                    //                                     .readdata
		input  wire        pulse_90deg_clk_clk,                         //                      pulse_90deg_clk.clk
		output wire [31:0] pulse_90deg_external_connection_export,      //      pulse_90deg_external_connection.export
		input  wire        pulse_90deg_reset_reset_n,                   //                    pulse_90deg_reset.reset_n
		input  wire [1:0]  pulse_90deg_s1_address,                      //                       pulse_90deg_s1.address
		input  wire        pulse_90deg_s1_write_n,                      //                                     .write_n
		input  wire [31:0] pulse_90deg_s1_writedata,                    //                                     .writedata
		input  wire        pulse_90deg_s1_chipselect,                   //                                     .chipselect
		output wire [31:0] pulse_90deg_s1_readdata,                     //                                     .readdata
		input  wire        pulse_t1_clk_clk,                            //                         pulse_t1_clk.clk
		output wire [31:0] pulse_t1_external_connection_export,         //         pulse_t1_external_connection.export
		input  wire        pulse_t1_reset_reset_n,                      //                       pulse_t1_reset.reset_n
		input  wire [1:0]  pulse_t1_s1_address,                         //                          pulse_t1_s1.address
		input  wire        pulse_t1_s1_write_n,                         //                                     .write_n
		input  wire [31:0] pulse_t1_s1_writedata,                       //                                     .writedata
		input  wire        pulse_t1_s1_chipselect,                      //                                     .chipselect
		output wire [31:0] pulse_t1_s1_readdata,                        //                                     .readdata
		input  wire        rx_delay_clk_clk,                            //                         rx_delay_clk.clk
		output wire [31:0] rx_delay_external_connection_export,         //         rx_delay_external_connection.export
		input  wire        rx_delay_reset_reset_n,                      //                       rx_delay_reset.reset_n
		input  wire [1:0]  rx_delay_s1_address,                         //                          rx_delay_s1.address
		input  wire        rx_delay_s1_write_n,                         //                                     .write_n
		input  wire [31:0] rx_delay_s1_writedata,                       //                                     .writedata
		input  wire        rx_delay_s1_chipselect,                      //                                     .chipselect
		output wire [31:0] rx_delay_s1_readdata,                        //                                     .readdata
		input  wire        samples_per_echo_clk_clk,                    //                 samples_per_echo_clk.clk
		output wire [31:0] samples_per_echo_external_connection_export, // samples_per_echo_external_connection.export
		input  wire        samples_per_echo_reset_reset_n,              //               samples_per_echo_reset.reset_n
		input  wire [1:0]  samples_per_echo_s1_address,                 //                  samples_per_echo_s1.address
		input  wire        samples_per_echo_s1_write_n,                 //                                     .write_n
		input  wire [31:0] samples_per_echo_s1_writedata,               //                                     .writedata
		input  wire        samples_per_echo_s1_chipselect,              //                                     .chipselect
		output wire [31:0] samples_per_echo_s1_readdata                 //                                     .readdata
	);

	soc_system_v5_nmr_parameters_adc_val_sub adc_val_sub (
		.clk        (adc_val_sub_clk_clk),                    //                 clk.clk
		.reset_n    (adc_val_sub_reset_reset_n),              //               reset.reset_n
		.address    (adc_val_sub_s1_address),                 //                  s1.address
		.write_n    (adc_val_sub_s1_write_n),                 //                    .write_n
		.writedata  (adc_val_sub_s1_writedata),               //                    .writedata
		.chipselect (adc_val_sub_s1_chipselect),              //                    .chipselect
		.readdata   (adc_val_sub_s1_readdata),                //                    .readdata
		.out_port   (adc_val_sub_external_connection_export)  // external_connection.export
	);

	soc_system_v5_nmr_parameters_delay_nosig delay_nosig (
		.clk        (delay_nosig_clk_clk),                    //                 clk.clk
		.reset_n    (delay_nosig_reset_reset_n),              //               reset.reset_n
		.address    (delay_nosig_s1_address),                 //                  s1.address
		.write_n    (delay_nosig_s1_write_n),                 //                    .write_n
		.writedata  (delay_nosig_s1_writedata),               //                    .writedata
		.chipselect (delay_nosig_s1_chipselect),              //                    .chipselect
		.readdata   (delay_nosig_s1_readdata),                //                    .readdata
		.out_port   (delay_nosig_external_connection_export)  // external_connection.export
	);

	soc_system_v5_nmr_parameters_delay_nosig delay_sig (
		.clk        (delay_sig_clk_clk),                    //                 clk.clk
		.reset_n    (delay_sig_reset_reset_n),              //               reset.reset_n
		.address    (delay_sig_s1_address),                 //                  s1.address
		.write_n    (delay_sig_s1_write_n),                 //                    .write_n
		.writedata  (delay_sig_s1_writedata),               //                    .writedata
		.chipselect (delay_sig_s1_chipselect),              //                    .chipselect
		.readdata   (delay_sig_s1_readdata),                //                    .readdata
		.out_port   (delay_sig_external_connection_export)  // external_connection.export
	);

	soc_system_v5_nmr_parameters_delay_t1 delay_t1 (
		.clk        (delay_t1_clk_clk),                    //                 clk.clk
		.reset_n    (delay_t1_reset_reset_n),              //               reset.reset_n
		.address    (delay_t1_s1_address),                 //                  s1.address
		.write_n    (delay_t1_s1_write_n),                 //                    .write_n
		.writedata  (delay_t1_s1_writedata),               //                    .writedata
		.chipselect (delay_t1_s1_chipselect),              //                    .chipselect
		.readdata   (delay_t1_s1_readdata),                //                    .readdata
		.out_port   (delay_t1_external_connection_export)  // external_connection.export
	);

	soc_system_v5_nmr_parameters_delay_t1 echoes_per_scan (
		.clk        (echoes_per_scan_clk_clk),                    //                 clk.clk
		.reset_n    (echoes_per_scan_reset_reset_n),              //               reset.reset_n
		.address    (echoes_per_scan_s1_address),                 //                  s1.address
		.write_n    (echoes_per_scan_s1_write_n),                 //                    .write_n
		.writedata  (echoes_per_scan_s1_writedata),               //                    .writedata
		.chipselect (echoes_per_scan_s1_chipselect),              //                    .chipselect
		.readdata   (echoes_per_scan_s1_readdata),                //                    .readdata
		.out_port   (echoes_per_scan_external_connection_export)  // external_connection.export
	);

	soc_system_v5_nmr_parameters_delay_t1 init_delay (
		.clk        (init_delay_clk_clk),                    //                 clk.clk
		.reset_n    (init_delay_reset_reset_n),              //               reset.reset_n
		.address    (init_delay_s1_address),                 //                  s1.address
		.write_n    (init_delay_s1_write_n),                 //                    .write_n
		.writedata  (init_delay_s1_writedata),               //                    .writedata
		.chipselect (init_delay_s1_chipselect),              //                    .chipselect
		.readdata   (init_delay_s1_readdata),                //                    .readdata
		.out_port   (init_delay_external_connection_export)  // external_connection.export
	);

	soc_system_v5_nmr_parameters_delay_nosig pulse_180deg (
		.clk        (pulse_180deg_clk_clk),                    //                 clk.clk
		.reset_n    (pulse_180deg_reset_reset_n),              //               reset.reset_n
		.address    (pulse_180deg_s1_address),                 //                  s1.address
		.write_n    (pulse_180deg_s1_write_n),                 //                    .write_n
		.writedata  (pulse_180deg_s1_writedata),               //                    .writedata
		.chipselect (pulse_180deg_s1_chipselect),              //                    .chipselect
		.readdata   (pulse_180deg_s1_readdata),                //                    .readdata
		.out_port   (pulse_180deg_external_connection_export)  // external_connection.export
	);

	soc_system_v5_nmr_parameters_delay_nosig pulse_90deg (
		.clk        (pulse_90deg_clk_clk),                    //                 clk.clk
		.reset_n    (pulse_90deg_reset_reset_n),              //               reset.reset_n
		.address    (pulse_90deg_s1_address),                 //                  s1.address
		.write_n    (pulse_90deg_s1_write_n),                 //                    .write_n
		.writedata  (pulse_90deg_s1_writedata),               //                    .writedata
		.chipselect (pulse_90deg_s1_chipselect),              //                    .chipselect
		.readdata   (pulse_90deg_s1_readdata),                //                    .readdata
		.out_port   (pulse_90deg_external_connection_export)  // external_connection.export
	);

	soc_system_v5_nmr_parameters_delay_t1 pulse_t1 (
		.clk        (pulse_t1_clk_clk),                    //                 clk.clk
		.reset_n    (pulse_t1_reset_reset_n),              //               reset.reset_n
		.address    (pulse_t1_s1_address),                 //                  s1.address
		.write_n    (pulse_t1_s1_write_n),                 //                    .write_n
		.writedata  (pulse_t1_s1_writedata),               //                    .writedata
		.chipselect (pulse_t1_s1_chipselect),              //                    .chipselect
		.readdata   (pulse_t1_s1_readdata),                //                    .readdata
		.out_port   (pulse_t1_external_connection_export)  // external_connection.export
	);

	soc_system_v5_nmr_parameters_delay_t1 rx_delay (
		.clk        (rx_delay_clk_clk),                    //                 clk.clk
		.reset_n    (rx_delay_reset_reset_n),              //               reset.reset_n
		.address    (rx_delay_s1_address),                 //                  s1.address
		.write_n    (rx_delay_s1_write_n),                 //                    .write_n
		.writedata  (rx_delay_s1_writedata),               //                    .writedata
		.chipselect (rx_delay_s1_chipselect),              //                    .chipselect
		.readdata   (rx_delay_s1_readdata),                //                    .readdata
		.out_port   (rx_delay_external_connection_export)  // external_connection.export
	);

	soc_system_v5_nmr_parameters_samples_per_echo samples_per_echo (
		.clk        (samples_per_echo_clk_clk),                    //                 clk.clk
		.reset_n    (samples_per_echo_reset_reset_n),              //               reset.reset_n
		.address    (samples_per_echo_s1_address),                 //                  s1.address
		.write_n    (samples_per_echo_s1_write_n),                 //                    .write_n
		.writedata  (samples_per_echo_s1_writedata),               //                    .writedata
		.chipselect (samples_per_echo_s1_chipselect),              //                    .chipselect
		.readdata   (samples_per_echo_s1_readdata),                //                    .readdata
		.out_port   (samples_per_echo_external_connection_export)  // external_connection.export
	);

endmodule
