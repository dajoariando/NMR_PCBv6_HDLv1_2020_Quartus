// FIR_filter_test_tb.v

// Generated using ACDS version 17.1 590

`timescale 1 ps / 1 ps
module FIR_filter_test_tb (
	);

	wire    fir_filter_test_inst_clk_bfm_clk_clk;       // FIR_filter_test_inst_clk_bfm:clk -> [FIR_filter_test_inst:clk_clk, FIR_filter_test_inst_reset_bfm:clk]
	wire    fir_filter_test_inst_reset_bfm_reset_reset; // FIR_filter_test_inst_reset_bfm:reset -> FIR_filter_test_inst:reset_reset_n

	FIR_filter_test fir_filter_test_inst (
		.clk_clk       (fir_filter_test_inst_clk_bfm_clk_clk),       //   clk.clk
		.reset_reset_n (fir_filter_test_inst_reset_bfm_reset_reset)  // reset.reset_n
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) fir_filter_test_inst_clk_bfm (
		.clk (fir_filter_test_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) fir_filter_test_inst_reset_bfm (
		.reset (fir_filter_test_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (fir_filter_test_inst_clk_bfm_clk_clk)        //   clk.clk
	);

endmodule
