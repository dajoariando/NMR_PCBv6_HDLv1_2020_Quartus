// system.v

// Generated using ACDS version 17.1 590

`timescale 1 ps / 1 ps
module system (
		input  wire        clk_clk,                 //                 clk.clk
		input  wire        dac_preamp_MISO,         //          dac_preamp.MISO
		output wire        dac_preamp_MOSI,         //                    .MOSI
		output wire        dac_preamp_SCLK,         //                    .SCLK
		output wire        dac_preamp_SS_n,         //                    .SS_n
		output wire [31:0] delay_nosig_export,      //         delay_nosig.export
		output wire [31:0] delay_sig_export,        //           delay_sig.export
		output wire [31:0] delay_t1_export,         //            delay_t1.export
		output wire [31:0] echoes_per_scan_export,  //     echoes_per_scan.export
		input  wire        i2c_ext_sda_in,          //             i2c_ext.sda_in
		input  wire        i2c_ext_scl_in,          //                    .scl_in
		output wire        i2c_ext_sda_oe,          //                    .sda_oe
		output wire        i2c_ext_scl_oe,          //                    .scl_oe
		input  wire        i2c_int_sda_in,          //             i2c_int.sda_in
		input  wire        i2c_int_scl_in,          //                    .scl_in
		output wire        i2c_int_sda_oe,          //                    .sda_oe
		output wire        i2c_int_scl_oe,          //                    .scl_oe
		output wire [31:0] init_delay_export,       //          init_delay.export
		output wire [0:0]  issp_source,             //                issp.source
		output wire [9:0]  led_export,              //                 led.export
		output wire        nmr_sys_pll_outclk0_clk, // nmr_sys_pll_outclk0.clk
		output wire [31:0] pulse_180deg_export,     //        pulse_180deg.export
		output wire [31:0] pulse_90deg_export,      //         pulse_90deg.export
		output wire [31:0] pulse_t1_export,         //            pulse_t1.export
		input  wire        reset_reset_n,           //               reset.reset_n
		output wire [31:0] samples_per_echo_export  //    samples_per_echo.export
	);

	wire  [63:0] nmr_sys_pll_reconfig_from_pll_reconfig_from_pll;                // nmr_sys_pll:reconfig_from_pll -> pll_reconfig_0:reconfig_from_pll
	wire  [63:0] pll_reconfig_0_reconfig_to_pll_reconfig_to_pll;                 // pll_reconfig_0:reconfig_to_pll -> nmr_sys_pll:reconfig_to_pll
	wire  [31:0] system_console_master_readdata;                                 // mm_interconnect_0:system_console_master_readdata -> system_console:master_readdata
	wire         system_console_master_waitrequest;                              // mm_interconnect_0:system_console_master_waitrequest -> system_console:master_waitrequest
	wire  [31:0] system_console_master_address;                                  // system_console:master_address -> mm_interconnect_0:system_console_master_address
	wire         system_console_master_read;                                     // system_console:master_read -> mm_interconnect_0:system_console_master_read
	wire   [3:0] system_console_master_byteenable;                               // system_console:master_byteenable -> mm_interconnect_0:system_console_master_byteenable
	wire         system_console_master_readdatavalid;                            // mm_interconnect_0:system_console_master_readdatavalid -> system_console:master_readdatavalid
	wire         system_console_master_write;                                    // system_console:master_write -> mm_interconnect_0:system_console_master_write
	wire  [31:0] system_console_master_writedata;                                // system_console:master_writedata -> mm_interconnect_0:system_console_master_writedata
	wire  [31:0] mm_interconnect_0_i2c_int_csr_readdata;                         // I2C_INT:readdata -> mm_interconnect_0:I2C_INT_csr_readdata
	wire   [3:0] mm_interconnect_0_i2c_int_csr_address;                          // mm_interconnect_0:I2C_INT_csr_address -> I2C_INT:addr
	wire         mm_interconnect_0_i2c_int_csr_read;                             // mm_interconnect_0:I2C_INT_csr_read -> I2C_INT:read
	wire         mm_interconnect_0_i2c_int_csr_write;                            // mm_interconnect_0:I2C_INT_csr_write -> I2C_INT:write
	wire  [31:0] mm_interconnect_0_i2c_int_csr_writedata;                        // mm_interconnect_0:I2C_INT_csr_writedata -> I2C_INT:writedata
	wire  [31:0] mm_interconnect_0_i2c_ext_csr_readdata;                         // I2C_EXT:readdata -> mm_interconnect_0:I2C_EXT_csr_readdata
	wire   [3:0] mm_interconnect_0_i2c_ext_csr_address;                          // mm_interconnect_0:I2C_EXT_csr_address -> I2C_EXT:addr
	wire         mm_interconnect_0_i2c_ext_csr_read;                             // mm_interconnect_0:I2C_EXT_csr_read -> I2C_EXT:read
	wire         mm_interconnect_0_i2c_ext_csr_write;                            // mm_interconnect_0:I2C_EXT_csr_write -> I2C_EXT:write
	wire  [31:0] mm_interconnect_0_i2c_ext_csr_writedata;                        // mm_interconnect_0:I2C_EXT_csr_writedata -> I2C_EXT:writedata
	wire         mm_interconnect_0_parameters_0_delay_nosig_s1_chipselect;       // mm_interconnect_0:parameters_0_delay_nosig_s1_chipselect -> parameters_0:delay_nosig_s1_chipselect
	wire  [31:0] mm_interconnect_0_parameters_0_delay_nosig_s1_readdata;         // parameters_0:delay_nosig_s1_readdata -> mm_interconnect_0:parameters_0_delay_nosig_s1_readdata
	wire   [1:0] mm_interconnect_0_parameters_0_delay_nosig_s1_address;          // mm_interconnect_0:parameters_0_delay_nosig_s1_address -> parameters_0:delay_nosig_s1_address
	wire         mm_interconnect_0_parameters_0_delay_nosig_s1_write;            // mm_interconnect_0:parameters_0_delay_nosig_s1_write -> parameters_0:delay_nosig_s1_write_n
	wire  [31:0] mm_interconnect_0_parameters_0_delay_nosig_s1_writedata;        // mm_interconnect_0:parameters_0_delay_nosig_s1_writedata -> parameters_0:delay_nosig_s1_writedata
	wire         mm_interconnect_0_parameters_0_delay_sig_s1_chipselect;         // mm_interconnect_0:parameters_0_delay_sig_s1_chipselect -> parameters_0:delay_sig_s1_chipselect
	wire  [31:0] mm_interconnect_0_parameters_0_delay_sig_s1_readdata;           // parameters_0:delay_sig_s1_readdata -> mm_interconnect_0:parameters_0_delay_sig_s1_readdata
	wire   [1:0] mm_interconnect_0_parameters_0_delay_sig_s1_address;            // mm_interconnect_0:parameters_0_delay_sig_s1_address -> parameters_0:delay_sig_s1_address
	wire         mm_interconnect_0_parameters_0_delay_sig_s1_write;              // mm_interconnect_0:parameters_0_delay_sig_s1_write -> parameters_0:delay_sig_s1_write_n
	wire  [31:0] mm_interconnect_0_parameters_0_delay_sig_s1_writedata;          // mm_interconnect_0:parameters_0_delay_sig_s1_writedata -> parameters_0:delay_sig_s1_writedata
	wire         mm_interconnect_0_parameters_0_delay_t1_s1_chipselect;          // mm_interconnect_0:parameters_0_delay_t1_s1_chipselect -> parameters_0:delay_t1_s1_chipselect
	wire  [31:0] mm_interconnect_0_parameters_0_delay_t1_s1_readdata;            // parameters_0:delay_t1_s1_readdata -> mm_interconnect_0:parameters_0_delay_t1_s1_readdata
	wire   [1:0] mm_interconnect_0_parameters_0_delay_t1_s1_address;             // mm_interconnect_0:parameters_0_delay_t1_s1_address -> parameters_0:delay_t1_s1_address
	wire         mm_interconnect_0_parameters_0_delay_t1_s1_write;               // mm_interconnect_0:parameters_0_delay_t1_s1_write -> parameters_0:delay_t1_s1_write_n
	wire  [31:0] mm_interconnect_0_parameters_0_delay_t1_s1_writedata;           // mm_interconnect_0:parameters_0_delay_t1_s1_writedata -> parameters_0:delay_t1_s1_writedata
	wire         mm_interconnect_0_parameters_0_echoes_per_scan_s1_chipselect;   // mm_interconnect_0:parameters_0_echoes_per_scan_s1_chipselect -> parameters_0:echoes_per_scan_s1_chipselect
	wire  [31:0] mm_interconnect_0_parameters_0_echoes_per_scan_s1_readdata;     // parameters_0:echoes_per_scan_s1_readdata -> mm_interconnect_0:parameters_0_echoes_per_scan_s1_readdata
	wire   [1:0] mm_interconnect_0_parameters_0_echoes_per_scan_s1_address;      // mm_interconnect_0:parameters_0_echoes_per_scan_s1_address -> parameters_0:echoes_per_scan_s1_address
	wire         mm_interconnect_0_parameters_0_echoes_per_scan_s1_write;        // mm_interconnect_0:parameters_0_echoes_per_scan_s1_write -> parameters_0:echoes_per_scan_s1_write_n
	wire  [31:0] mm_interconnect_0_parameters_0_echoes_per_scan_s1_writedata;    // mm_interconnect_0:parameters_0_echoes_per_scan_s1_writedata -> parameters_0:echoes_per_scan_s1_writedata
	wire         mm_interconnect_0_parameters_0_init_delay_s1_chipselect;        // mm_interconnect_0:parameters_0_init_delay_s1_chipselect -> parameters_0:init_delay_s1_chipselect
	wire  [31:0] mm_interconnect_0_parameters_0_init_delay_s1_readdata;          // parameters_0:init_delay_s1_readdata -> mm_interconnect_0:parameters_0_init_delay_s1_readdata
	wire   [1:0] mm_interconnect_0_parameters_0_init_delay_s1_address;           // mm_interconnect_0:parameters_0_init_delay_s1_address -> parameters_0:init_delay_s1_address
	wire         mm_interconnect_0_parameters_0_init_delay_s1_write;             // mm_interconnect_0:parameters_0_init_delay_s1_write -> parameters_0:init_delay_s1_write_n
	wire  [31:0] mm_interconnect_0_parameters_0_init_delay_s1_writedata;         // mm_interconnect_0:parameters_0_init_delay_s1_writedata -> parameters_0:init_delay_s1_writedata
	wire  [31:0] mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_readdata;    // pll_reconfig_0:mgmt_readdata -> mm_interconnect_0:pll_reconfig_0_mgmt_avalon_slave_readdata
	wire         mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_waitrequest; // pll_reconfig_0:mgmt_waitrequest -> mm_interconnect_0:pll_reconfig_0_mgmt_avalon_slave_waitrequest
	wire   [5:0] mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_address;     // mm_interconnect_0:pll_reconfig_0_mgmt_avalon_slave_address -> pll_reconfig_0:mgmt_address
	wire         mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_read;        // mm_interconnect_0:pll_reconfig_0_mgmt_avalon_slave_read -> pll_reconfig_0:mgmt_read
	wire         mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_write;       // mm_interconnect_0:pll_reconfig_0_mgmt_avalon_slave_write -> pll_reconfig_0:mgmt_write
	wire  [31:0] mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_writedata;   // mm_interconnect_0:pll_reconfig_0_mgmt_avalon_slave_writedata -> pll_reconfig_0:mgmt_writedata
	wire         mm_interconnect_0_parameters_0_pulse_180deg_s1_chipselect;      // mm_interconnect_0:parameters_0_pulse_180deg_s1_chipselect -> parameters_0:pulse_180deg_s1_chipselect
	wire  [31:0] mm_interconnect_0_parameters_0_pulse_180deg_s1_readdata;        // parameters_0:pulse_180deg_s1_readdata -> mm_interconnect_0:parameters_0_pulse_180deg_s1_readdata
	wire   [1:0] mm_interconnect_0_parameters_0_pulse_180deg_s1_address;         // mm_interconnect_0:parameters_0_pulse_180deg_s1_address -> parameters_0:pulse_180deg_s1_address
	wire         mm_interconnect_0_parameters_0_pulse_180deg_s1_write;           // mm_interconnect_0:parameters_0_pulse_180deg_s1_write -> parameters_0:pulse_180deg_s1_write_n
	wire  [31:0] mm_interconnect_0_parameters_0_pulse_180deg_s1_writedata;       // mm_interconnect_0:parameters_0_pulse_180deg_s1_writedata -> parameters_0:pulse_180deg_s1_writedata
	wire         mm_interconnect_0_parameters_0_pulse_90deg_s1_chipselect;       // mm_interconnect_0:parameters_0_pulse_90deg_s1_chipselect -> parameters_0:pulse_90deg_s1_chipselect
	wire  [31:0] mm_interconnect_0_parameters_0_pulse_90deg_s1_readdata;         // parameters_0:pulse_90deg_s1_readdata -> mm_interconnect_0:parameters_0_pulse_90deg_s1_readdata
	wire   [1:0] mm_interconnect_0_parameters_0_pulse_90deg_s1_address;          // mm_interconnect_0:parameters_0_pulse_90deg_s1_address -> parameters_0:pulse_90deg_s1_address
	wire         mm_interconnect_0_parameters_0_pulse_90deg_s1_write;            // mm_interconnect_0:parameters_0_pulse_90deg_s1_write -> parameters_0:pulse_90deg_s1_write_n
	wire  [31:0] mm_interconnect_0_parameters_0_pulse_90deg_s1_writedata;        // mm_interconnect_0:parameters_0_pulse_90deg_s1_writedata -> parameters_0:pulse_90deg_s1_writedata
	wire         mm_interconnect_0_parameters_0_pulse_t1_s1_chipselect;          // mm_interconnect_0:parameters_0_pulse_t1_s1_chipselect -> parameters_0:pulse_t1_s1_chipselect
	wire  [31:0] mm_interconnect_0_parameters_0_pulse_t1_s1_readdata;            // parameters_0:pulse_t1_s1_readdata -> mm_interconnect_0:parameters_0_pulse_t1_s1_readdata
	wire   [1:0] mm_interconnect_0_parameters_0_pulse_t1_s1_address;             // mm_interconnect_0:parameters_0_pulse_t1_s1_address -> parameters_0:pulse_t1_s1_address
	wire         mm_interconnect_0_parameters_0_pulse_t1_s1_write;               // mm_interconnect_0:parameters_0_pulse_t1_s1_write -> parameters_0:pulse_t1_s1_write_n
	wire  [31:0] mm_interconnect_0_parameters_0_pulse_t1_s1_writedata;           // mm_interconnect_0:parameters_0_pulse_t1_s1_writedata -> parameters_0:pulse_t1_s1_writedata
	wire         mm_interconnect_0_led_s1_chipselect;                            // mm_interconnect_0:led_s1_chipselect -> led:chipselect
	wire  [31:0] mm_interconnect_0_led_s1_readdata;                              // led:readdata -> mm_interconnect_0:led_s1_readdata
	wire   [1:0] mm_interconnect_0_led_s1_address;                               // mm_interconnect_0:led_s1_address -> led:address
	wire         mm_interconnect_0_led_s1_write;                                 // mm_interconnect_0:led_s1_write -> led:write_n
	wire  [31:0] mm_interconnect_0_led_s1_writedata;                             // mm_interconnect_0:led_s1_writedata -> led:writedata
	wire         mm_interconnect_0_parameters_0_samples_per_echo_s1_chipselect;  // mm_interconnect_0:parameters_0_samples_per_echo_s1_chipselect -> parameters_0:samples_per_echo_s1_chipselect
	wire  [31:0] mm_interconnect_0_parameters_0_samples_per_echo_s1_readdata;    // parameters_0:samples_per_echo_s1_readdata -> mm_interconnect_0:parameters_0_samples_per_echo_s1_readdata
	wire   [1:0] mm_interconnect_0_parameters_0_samples_per_echo_s1_address;     // mm_interconnect_0:parameters_0_samples_per_echo_s1_address -> parameters_0:samples_per_echo_s1_address
	wire         mm_interconnect_0_parameters_0_samples_per_echo_s1_write;       // mm_interconnect_0:parameters_0_samples_per_echo_s1_write -> parameters_0:samples_per_echo_s1_write_n
	wire  [31:0] mm_interconnect_0_parameters_0_samples_per_echo_s1_writedata;   // mm_interconnect_0:parameters_0_samples_per_echo_s1_writedata -> parameters_0:samples_per_echo_s1_writedata
	wire         mm_interconnect_0_dac_preamp_spi_control_port_chipselect;       // mm_interconnect_0:dac_preamp_spi_control_port_chipselect -> dac_preamp:spi_select
	wire  [31:0] mm_interconnect_0_dac_preamp_spi_control_port_readdata;         // dac_preamp:data_to_cpu -> mm_interconnect_0:dac_preamp_spi_control_port_readdata
	wire   [2:0] mm_interconnect_0_dac_preamp_spi_control_port_address;          // mm_interconnect_0:dac_preamp_spi_control_port_address -> dac_preamp:mem_addr
	wire         mm_interconnect_0_dac_preamp_spi_control_port_read;             // mm_interconnect_0:dac_preamp_spi_control_port_read -> dac_preamp:read_n
	wire         mm_interconnect_0_dac_preamp_spi_control_port_write;            // mm_interconnect_0:dac_preamp_spi_control_port_write -> dac_preamp:write_n
	wire  [31:0] mm_interconnect_0_dac_preamp_spi_control_port_writedata;        // mm_interconnect_0:dac_preamp_spi_control_port_writedata -> dac_preamp:data_from_cpu
	wire         rst_controller_reset_out_reset;                                 // rst_controller:reset_out -> [I2C_EXT:rst_n, I2C_INT:rst_n, dac_preamp:reset_n, led:reset_n, mm_interconnect_0:I2C_INT_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_0:system_console_clk_reset_reset_bridge_in_reset_reset, pll_reconfig_0:mgmt_reset]

	altera_avalon_i2c #(
		.USE_AV_ST       (0),
		.FIFO_DEPTH      (16),
		.FIFO_DEPTH_LOG2 (4)
	) i2c_ext (
		.clk       (clk_clk),                                 //            clock.clk
		.rst_n     (~rst_controller_reset_out_reset),         //       reset_sink.reset_n
		.intr      (),                                        // interrupt_sender.irq
		.addr      (mm_interconnect_0_i2c_ext_csr_address),   //              csr.address
		.read      (mm_interconnect_0_i2c_ext_csr_read),      //                 .read
		.write     (mm_interconnect_0_i2c_ext_csr_write),     //                 .write
		.writedata (mm_interconnect_0_i2c_ext_csr_writedata), //                 .writedata
		.readdata  (mm_interconnect_0_i2c_ext_csr_readdata),  //                 .readdata
		.sda_in    (i2c_ext_sda_in),                          //       i2c_serial.sda_in
		.scl_in    (i2c_ext_scl_in),                          //                 .scl_in
		.sda_oe    (i2c_ext_sda_oe),                          //                 .sda_oe
		.scl_oe    (i2c_ext_scl_oe),                          //                 .scl_oe
		.src_data  (),                                        //      (terminated)
		.src_valid (),                                        //      (terminated)
		.src_ready (1'b0),                                    //      (terminated)
		.snk_data  (16'b0000000000000000),                    //      (terminated)
		.snk_valid (1'b0),                                    //      (terminated)
		.snk_ready ()                                         //      (terminated)
	);

	altera_avalon_i2c #(
		.USE_AV_ST       (0),
		.FIFO_DEPTH      (16),
		.FIFO_DEPTH_LOG2 (4)
	) i2c_int (
		.clk       (clk_clk),                                 //            clock.clk
		.rst_n     (~rst_controller_reset_out_reset),         //       reset_sink.reset_n
		.intr      (),                                        // interrupt_sender.irq
		.addr      (mm_interconnect_0_i2c_int_csr_address),   //              csr.address
		.read      (mm_interconnect_0_i2c_int_csr_read),      //                 .read
		.write     (mm_interconnect_0_i2c_int_csr_write),     //                 .write
		.writedata (mm_interconnect_0_i2c_int_csr_writedata), //                 .writedata
		.readdata  (mm_interconnect_0_i2c_int_csr_readdata),  //                 .readdata
		.sda_in    (i2c_int_sda_in),                          //       i2c_serial.sda_in
		.scl_in    (i2c_int_scl_in),                          //                 .scl_in
		.sda_oe    (i2c_int_sda_oe),                          //                 .sda_oe
		.scl_oe    (i2c_int_scl_oe),                          //                 .scl_oe
		.src_data  (),                                        //      (terminated)
		.src_valid (),                                        //      (terminated)
		.src_ready (1'b0),                                    //      (terminated)
		.snk_data  (16'b0000000000000000),                    //      (terminated)
		.snk_valid (1'b0),                                    //      (terminated)
		.snk_ready ()                                         //      (terminated)
	);

	system_dac_preamp dac_preamp (
		.clk           (clk_clk),                                                  //              clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                          //            reset.reset_n
		.data_from_cpu (mm_interconnect_0_dac_preamp_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_0_dac_preamp_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_0_dac_preamp_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_0_dac_preamp_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_0_dac_preamp_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_0_dac_preamp_spi_control_port_write),     //                 .write_n
		.irq           (),                                                         //              irq.irq
		.MISO          (dac_preamp_MISO),                                          //         external.export
		.MOSI          (dac_preamp_MOSI),                                          //                 .export
		.SCLK          (dac_preamp_SCLK),                                          //                 .export
		.SS_n          (dac_preamp_SS_n)                                           //                 .export
	);

	altsource_probe_top #(
		.sld_auto_instance_index ("YES"),
		.sld_instance_index      (0),
		.instance_id             ("NONE"),
		.probe_width             (0),
		.source_width            (1),
		.source_initial_value    ("0"),
		.enable_metastability    ("NO")
	) in_system_sources_probes_0 (
		.source     (issp_source), // sources.source
		.source_ena (1'b1)         // (terminated)
	);

	system_led led (
		.clk        (clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_s1_readdata),   //                    .readdata
		.out_port   (led_export)                           // external_connection.export
	);

	system_nmr_sys_pll nmr_sys_pll (
		.refclk            (clk_clk),                                         //            refclk.clk
		.rst               (~reset_reset_n),                                  //             reset.reset
		.outclk_0          (nmr_sys_pll_outclk0_clk),                         //           outclk0.clk
		.reconfig_to_pll   (pll_reconfig_0_reconfig_to_pll_reconfig_to_pll),  //   reconfig_to_pll.reconfig_to_pll
		.reconfig_from_pll (nmr_sys_pll_reconfig_from_pll_reconfig_from_pll), // reconfig_from_pll.reconfig_from_pll
		.locked            ()                                                 //       (terminated)
	);

	system_parameters_0 parameters_0 (
		.clk_clk                                     (clk_clk),                                                       //                                  clk.clk
		.delay_nosig_external_connection_export      (delay_nosig_export),                                            //      delay_nosig_external_connection.export
		.delay_nosig_s1_address                      (mm_interconnect_0_parameters_0_delay_nosig_s1_address),         //                       delay_nosig_s1.address
		.delay_nosig_s1_write_n                      (~mm_interconnect_0_parameters_0_delay_nosig_s1_write),          //                                     .write_n
		.delay_nosig_s1_writedata                    (mm_interconnect_0_parameters_0_delay_nosig_s1_writedata),       //                                     .writedata
		.delay_nosig_s1_chipselect                   (mm_interconnect_0_parameters_0_delay_nosig_s1_chipselect),      //                                     .chipselect
		.delay_nosig_s1_readdata                     (mm_interconnect_0_parameters_0_delay_nosig_s1_readdata),        //                                     .readdata
		.delay_sig_external_connection_export        (delay_sig_export),                                              //        delay_sig_external_connection.export
		.delay_sig_s1_address                        (mm_interconnect_0_parameters_0_delay_sig_s1_address),           //                         delay_sig_s1.address
		.delay_sig_s1_write_n                        (~mm_interconnect_0_parameters_0_delay_sig_s1_write),            //                                     .write_n
		.delay_sig_s1_writedata                      (mm_interconnect_0_parameters_0_delay_sig_s1_writedata),         //                                     .writedata
		.delay_sig_s1_chipselect                     (mm_interconnect_0_parameters_0_delay_sig_s1_chipselect),        //                                     .chipselect
		.delay_sig_s1_readdata                       (mm_interconnect_0_parameters_0_delay_sig_s1_readdata),          //                                     .readdata
		.delay_t1_external_connection_export         (delay_t1_export),                                               //         delay_t1_external_connection.export
		.delay_t1_s1_address                         (mm_interconnect_0_parameters_0_delay_t1_s1_address),            //                          delay_t1_s1.address
		.delay_t1_s1_write_n                         (~mm_interconnect_0_parameters_0_delay_t1_s1_write),             //                                     .write_n
		.delay_t1_s1_writedata                       (mm_interconnect_0_parameters_0_delay_t1_s1_writedata),          //                                     .writedata
		.delay_t1_s1_chipselect                      (mm_interconnect_0_parameters_0_delay_t1_s1_chipselect),         //                                     .chipselect
		.delay_t1_s1_readdata                        (mm_interconnect_0_parameters_0_delay_t1_s1_readdata),           //                                     .readdata
		.echoes_per_scan_external_connection_export  (echoes_per_scan_export),                                        //  echoes_per_scan_external_connection.export
		.echoes_per_scan_s1_address                  (mm_interconnect_0_parameters_0_echoes_per_scan_s1_address),     //                   echoes_per_scan_s1.address
		.echoes_per_scan_s1_write_n                  (~mm_interconnect_0_parameters_0_echoes_per_scan_s1_write),      //                                     .write_n
		.echoes_per_scan_s1_writedata                (mm_interconnect_0_parameters_0_echoes_per_scan_s1_writedata),   //                                     .writedata
		.echoes_per_scan_s1_chipselect               (mm_interconnect_0_parameters_0_echoes_per_scan_s1_chipselect),  //                                     .chipselect
		.echoes_per_scan_s1_readdata                 (mm_interconnect_0_parameters_0_echoes_per_scan_s1_readdata),    //                                     .readdata
		.init_delay_external_connection_export       (init_delay_export),                                             //       init_delay_external_connection.export
		.init_delay_s1_address                       (mm_interconnect_0_parameters_0_init_delay_s1_address),          //                        init_delay_s1.address
		.init_delay_s1_write_n                       (~mm_interconnect_0_parameters_0_init_delay_s1_write),           //                                     .write_n
		.init_delay_s1_writedata                     (mm_interconnect_0_parameters_0_init_delay_s1_writedata),        //                                     .writedata
		.init_delay_s1_chipselect                    (mm_interconnect_0_parameters_0_init_delay_s1_chipselect),       //                                     .chipselect
		.init_delay_s1_readdata                      (mm_interconnect_0_parameters_0_init_delay_s1_readdata),         //                                     .readdata
		.pulse_180deg_external_connection_export     (pulse_180deg_export),                                           //     pulse_180deg_external_connection.export
		.pulse_180deg_s1_address                     (mm_interconnect_0_parameters_0_pulse_180deg_s1_address),        //                      pulse_180deg_s1.address
		.pulse_180deg_s1_write_n                     (~mm_interconnect_0_parameters_0_pulse_180deg_s1_write),         //                                     .write_n
		.pulse_180deg_s1_writedata                   (mm_interconnect_0_parameters_0_pulse_180deg_s1_writedata),      //                                     .writedata
		.pulse_180deg_s1_chipselect                  (mm_interconnect_0_parameters_0_pulse_180deg_s1_chipselect),     //                                     .chipselect
		.pulse_180deg_s1_readdata                    (mm_interconnect_0_parameters_0_pulse_180deg_s1_readdata),       //                                     .readdata
		.pulse_90deg_external_connection_export      (pulse_90deg_export),                                            //      pulse_90deg_external_connection.export
		.pulse_90deg_s1_address                      (mm_interconnect_0_parameters_0_pulse_90deg_s1_address),         //                       pulse_90deg_s1.address
		.pulse_90deg_s1_write_n                      (~mm_interconnect_0_parameters_0_pulse_90deg_s1_write),          //                                     .write_n
		.pulse_90deg_s1_writedata                    (mm_interconnect_0_parameters_0_pulse_90deg_s1_writedata),       //                                     .writedata
		.pulse_90deg_s1_chipselect                   (mm_interconnect_0_parameters_0_pulse_90deg_s1_chipselect),      //                                     .chipselect
		.pulse_90deg_s1_readdata                     (mm_interconnect_0_parameters_0_pulse_90deg_s1_readdata),        //                                     .readdata
		.pulse_t1_external_connection_export         (pulse_t1_export),                                               //         pulse_t1_external_connection.export
		.pulse_t1_s1_address                         (mm_interconnect_0_parameters_0_pulse_t1_s1_address),            //                          pulse_t1_s1.address
		.pulse_t1_s1_write_n                         (~mm_interconnect_0_parameters_0_pulse_t1_s1_write),             //                                     .write_n
		.pulse_t1_s1_writedata                       (mm_interconnect_0_parameters_0_pulse_t1_s1_writedata),          //                                     .writedata
		.pulse_t1_s1_chipselect                      (mm_interconnect_0_parameters_0_pulse_t1_s1_chipselect),         //                                     .chipselect
		.pulse_t1_s1_readdata                        (mm_interconnect_0_parameters_0_pulse_t1_s1_readdata),           //                                     .readdata
		.reset_reset_n                               (reset_reset_n),                                                 //                                reset.reset_n
		.samples_per_echo_external_connection_export (samples_per_echo_export),                                       // samples_per_echo_external_connection.export
		.samples_per_echo_s1_address                 (mm_interconnect_0_parameters_0_samples_per_echo_s1_address),    //                  samples_per_echo_s1.address
		.samples_per_echo_s1_write_n                 (~mm_interconnect_0_parameters_0_samples_per_echo_s1_write),     //                                     .write_n
		.samples_per_echo_s1_writedata               (mm_interconnect_0_parameters_0_samples_per_echo_s1_writedata),  //                                     .writedata
		.samples_per_echo_s1_chipselect              (mm_interconnect_0_parameters_0_samples_per_echo_s1_chipselect), //                                     .chipselect
		.samples_per_echo_s1_readdata                (mm_interconnect_0_parameters_0_samples_per_echo_s1_readdata)    //                                     .readdata
	);

	altera_pll_reconfig_top #(
		.device_family       ("Cyclone V"),
		.ENABLE_MIF          (0),
		.MIF_FILE_NAME       (""),
		.ENABLE_BYTEENABLE   (0),
		.BYTEENABLE_WIDTH    (4),
		.RECONFIG_ADDR_WIDTH (6),
		.RECONFIG_DATA_WIDTH (32),
		.reconf_width        (64),
		.WAIT_FOR_LOCK       (1)
	) pll_reconfig_0 (
		.mgmt_clk          (clk_clk),                                                        //          mgmt_clk.clk
		.mgmt_reset        (rst_controller_reset_out_reset),                                 //        mgmt_reset.reset
		.mgmt_waitrequest  (mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_waitrequest), // mgmt_avalon_slave.waitrequest
		.mgmt_read         (mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_read),        //                  .read
		.mgmt_write        (mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_write),       //                  .write
		.mgmt_readdata     (mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_readdata),    //                  .readdata
		.mgmt_address      (mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_address),     //                  .address
		.mgmt_writedata    (mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_writedata),   //                  .writedata
		.reconfig_to_pll   (pll_reconfig_0_reconfig_to_pll_reconfig_to_pll),                 //   reconfig_to_pll.reconfig_to_pll
		.reconfig_from_pll (nmr_sys_pll_reconfig_from_pll_reconfig_from_pll),                // reconfig_from_pll.reconfig_from_pll
		.mgmt_byteenable   (4'b0000)                                                         //       (terminated)
	);

	system_system_console #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) system_console (
		.clk_clk              (clk_clk),                             //          clk.clk
		.clk_reset_reset      (~reset_reset_n),                      //    clk_reset.reset
		.master_address       (system_console_master_address),       //       master.address
		.master_readdata      (system_console_master_readdata),      //             .readdata
		.master_read          (system_console_master_read),          //             .read
		.master_write         (system_console_master_write),         //             .write
		.master_writedata     (system_console_master_writedata),     //             .writedata
		.master_waitrequest   (system_console_master_waitrequest),   //             .waitrequest
		.master_readdatavalid (system_console_master_readdatavalid), //             .readdatavalid
		.master_byteenable    (system_console_master_byteenable),    //             .byteenable
		.master_reset_reset   ()                                     // master_reset.reset
	);

	system_mm_interconnect_0 mm_interconnect_0 (
		.clk_in_clk_clk                                       (clk_clk),                                                        //                                     clk_in_clk.clk
		.I2C_INT_reset_sink_reset_bridge_in_reset_reset       (rst_controller_reset_out_reset),                                 //       I2C_INT_reset_sink_reset_bridge_in_reset.reset
		.system_console_clk_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                 // system_console_clk_reset_reset_bridge_in_reset.reset
		.system_console_master_address                        (system_console_master_address),                                  //                          system_console_master.address
		.system_console_master_waitrequest                    (system_console_master_waitrequest),                              //                                               .waitrequest
		.system_console_master_byteenable                     (system_console_master_byteenable),                               //                                               .byteenable
		.system_console_master_read                           (system_console_master_read),                                     //                                               .read
		.system_console_master_readdata                       (system_console_master_readdata),                                 //                                               .readdata
		.system_console_master_readdatavalid                  (system_console_master_readdatavalid),                            //                                               .readdatavalid
		.system_console_master_write                          (system_console_master_write),                                    //                                               .write
		.system_console_master_writedata                      (system_console_master_writedata),                                //                                               .writedata
		.dac_preamp_spi_control_port_address                  (mm_interconnect_0_dac_preamp_spi_control_port_address),          //                    dac_preamp_spi_control_port.address
		.dac_preamp_spi_control_port_write                    (mm_interconnect_0_dac_preamp_spi_control_port_write),            //                                               .write
		.dac_preamp_spi_control_port_read                     (mm_interconnect_0_dac_preamp_spi_control_port_read),             //                                               .read
		.dac_preamp_spi_control_port_readdata                 (mm_interconnect_0_dac_preamp_spi_control_port_readdata),         //                                               .readdata
		.dac_preamp_spi_control_port_writedata                (mm_interconnect_0_dac_preamp_spi_control_port_writedata),        //                                               .writedata
		.dac_preamp_spi_control_port_chipselect               (mm_interconnect_0_dac_preamp_spi_control_port_chipselect),       //                                               .chipselect
		.I2C_EXT_csr_address                                  (mm_interconnect_0_i2c_ext_csr_address),                          //                                    I2C_EXT_csr.address
		.I2C_EXT_csr_write                                    (mm_interconnect_0_i2c_ext_csr_write),                            //                                               .write
		.I2C_EXT_csr_read                                     (mm_interconnect_0_i2c_ext_csr_read),                             //                                               .read
		.I2C_EXT_csr_readdata                                 (mm_interconnect_0_i2c_ext_csr_readdata),                         //                                               .readdata
		.I2C_EXT_csr_writedata                                (mm_interconnect_0_i2c_ext_csr_writedata),                        //                                               .writedata
		.I2C_INT_csr_address                                  (mm_interconnect_0_i2c_int_csr_address),                          //                                    I2C_INT_csr.address
		.I2C_INT_csr_write                                    (mm_interconnect_0_i2c_int_csr_write),                            //                                               .write
		.I2C_INT_csr_read                                     (mm_interconnect_0_i2c_int_csr_read),                             //                                               .read
		.I2C_INT_csr_readdata                                 (mm_interconnect_0_i2c_int_csr_readdata),                         //                                               .readdata
		.I2C_INT_csr_writedata                                (mm_interconnect_0_i2c_int_csr_writedata),                        //                                               .writedata
		.led_s1_address                                       (mm_interconnect_0_led_s1_address),                               //                                         led_s1.address
		.led_s1_write                                         (mm_interconnect_0_led_s1_write),                                 //                                               .write
		.led_s1_readdata                                      (mm_interconnect_0_led_s1_readdata),                              //                                               .readdata
		.led_s1_writedata                                     (mm_interconnect_0_led_s1_writedata),                             //                                               .writedata
		.led_s1_chipselect                                    (mm_interconnect_0_led_s1_chipselect),                            //                                               .chipselect
		.parameters_0_delay_nosig_s1_address                  (mm_interconnect_0_parameters_0_delay_nosig_s1_address),          //                    parameters_0_delay_nosig_s1.address
		.parameters_0_delay_nosig_s1_write                    (mm_interconnect_0_parameters_0_delay_nosig_s1_write),            //                                               .write
		.parameters_0_delay_nosig_s1_readdata                 (mm_interconnect_0_parameters_0_delay_nosig_s1_readdata),         //                                               .readdata
		.parameters_0_delay_nosig_s1_writedata                (mm_interconnect_0_parameters_0_delay_nosig_s1_writedata),        //                                               .writedata
		.parameters_0_delay_nosig_s1_chipselect               (mm_interconnect_0_parameters_0_delay_nosig_s1_chipselect),       //                                               .chipselect
		.parameters_0_delay_sig_s1_address                    (mm_interconnect_0_parameters_0_delay_sig_s1_address),            //                      parameters_0_delay_sig_s1.address
		.parameters_0_delay_sig_s1_write                      (mm_interconnect_0_parameters_0_delay_sig_s1_write),              //                                               .write
		.parameters_0_delay_sig_s1_readdata                   (mm_interconnect_0_parameters_0_delay_sig_s1_readdata),           //                                               .readdata
		.parameters_0_delay_sig_s1_writedata                  (mm_interconnect_0_parameters_0_delay_sig_s1_writedata),          //                                               .writedata
		.parameters_0_delay_sig_s1_chipselect                 (mm_interconnect_0_parameters_0_delay_sig_s1_chipselect),         //                                               .chipselect
		.parameters_0_delay_t1_s1_address                     (mm_interconnect_0_parameters_0_delay_t1_s1_address),             //                       parameters_0_delay_t1_s1.address
		.parameters_0_delay_t1_s1_write                       (mm_interconnect_0_parameters_0_delay_t1_s1_write),               //                                               .write
		.parameters_0_delay_t1_s1_readdata                    (mm_interconnect_0_parameters_0_delay_t1_s1_readdata),            //                                               .readdata
		.parameters_0_delay_t1_s1_writedata                   (mm_interconnect_0_parameters_0_delay_t1_s1_writedata),           //                                               .writedata
		.parameters_0_delay_t1_s1_chipselect                  (mm_interconnect_0_parameters_0_delay_t1_s1_chipselect),          //                                               .chipselect
		.parameters_0_echoes_per_scan_s1_address              (mm_interconnect_0_parameters_0_echoes_per_scan_s1_address),      //                parameters_0_echoes_per_scan_s1.address
		.parameters_0_echoes_per_scan_s1_write                (mm_interconnect_0_parameters_0_echoes_per_scan_s1_write),        //                                               .write
		.parameters_0_echoes_per_scan_s1_readdata             (mm_interconnect_0_parameters_0_echoes_per_scan_s1_readdata),     //                                               .readdata
		.parameters_0_echoes_per_scan_s1_writedata            (mm_interconnect_0_parameters_0_echoes_per_scan_s1_writedata),    //                                               .writedata
		.parameters_0_echoes_per_scan_s1_chipselect           (mm_interconnect_0_parameters_0_echoes_per_scan_s1_chipselect),   //                                               .chipselect
		.parameters_0_init_delay_s1_address                   (mm_interconnect_0_parameters_0_init_delay_s1_address),           //                     parameters_0_init_delay_s1.address
		.parameters_0_init_delay_s1_write                     (mm_interconnect_0_parameters_0_init_delay_s1_write),             //                                               .write
		.parameters_0_init_delay_s1_readdata                  (mm_interconnect_0_parameters_0_init_delay_s1_readdata),          //                                               .readdata
		.parameters_0_init_delay_s1_writedata                 (mm_interconnect_0_parameters_0_init_delay_s1_writedata),         //                                               .writedata
		.parameters_0_init_delay_s1_chipselect                (mm_interconnect_0_parameters_0_init_delay_s1_chipselect),        //                                               .chipselect
		.parameters_0_pulse_180deg_s1_address                 (mm_interconnect_0_parameters_0_pulse_180deg_s1_address),         //                   parameters_0_pulse_180deg_s1.address
		.parameters_0_pulse_180deg_s1_write                   (mm_interconnect_0_parameters_0_pulse_180deg_s1_write),           //                                               .write
		.parameters_0_pulse_180deg_s1_readdata                (mm_interconnect_0_parameters_0_pulse_180deg_s1_readdata),        //                                               .readdata
		.parameters_0_pulse_180deg_s1_writedata               (mm_interconnect_0_parameters_0_pulse_180deg_s1_writedata),       //                                               .writedata
		.parameters_0_pulse_180deg_s1_chipselect              (mm_interconnect_0_parameters_0_pulse_180deg_s1_chipselect),      //                                               .chipselect
		.parameters_0_pulse_90deg_s1_address                  (mm_interconnect_0_parameters_0_pulse_90deg_s1_address),          //                    parameters_0_pulse_90deg_s1.address
		.parameters_0_pulse_90deg_s1_write                    (mm_interconnect_0_parameters_0_pulse_90deg_s1_write),            //                                               .write
		.parameters_0_pulse_90deg_s1_readdata                 (mm_interconnect_0_parameters_0_pulse_90deg_s1_readdata),         //                                               .readdata
		.parameters_0_pulse_90deg_s1_writedata                (mm_interconnect_0_parameters_0_pulse_90deg_s1_writedata),        //                                               .writedata
		.parameters_0_pulse_90deg_s1_chipselect               (mm_interconnect_0_parameters_0_pulse_90deg_s1_chipselect),       //                                               .chipselect
		.parameters_0_pulse_t1_s1_address                     (mm_interconnect_0_parameters_0_pulse_t1_s1_address),             //                       parameters_0_pulse_t1_s1.address
		.parameters_0_pulse_t1_s1_write                       (mm_interconnect_0_parameters_0_pulse_t1_s1_write),               //                                               .write
		.parameters_0_pulse_t1_s1_readdata                    (mm_interconnect_0_parameters_0_pulse_t1_s1_readdata),            //                                               .readdata
		.parameters_0_pulse_t1_s1_writedata                   (mm_interconnect_0_parameters_0_pulse_t1_s1_writedata),           //                                               .writedata
		.parameters_0_pulse_t1_s1_chipselect                  (mm_interconnect_0_parameters_0_pulse_t1_s1_chipselect),          //                                               .chipselect
		.parameters_0_samples_per_echo_s1_address             (mm_interconnect_0_parameters_0_samples_per_echo_s1_address),     //               parameters_0_samples_per_echo_s1.address
		.parameters_0_samples_per_echo_s1_write               (mm_interconnect_0_parameters_0_samples_per_echo_s1_write),       //                                               .write
		.parameters_0_samples_per_echo_s1_readdata            (mm_interconnect_0_parameters_0_samples_per_echo_s1_readdata),    //                                               .readdata
		.parameters_0_samples_per_echo_s1_writedata           (mm_interconnect_0_parameters_0_samples_per_echo_s1_writedata),   //                                               .writedata
		.parameters_0_samples_per_echo_s1_chipselect          (mm_interconnect_0_parameters_0_samples_per_echo_s1_chipselect),  //                                               .chipselect
		.pll_reconfig_0_mgmt_avalon_slave_address             (mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_address),     //               pll_reconfig_0_mgmt_avalon_slave.address
		.pll_reconfig_0_mgmt_avalon_slave_write               (mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_write),       //                                               .write
		.pll_reconfig_0_mgmt_avalon_slave_read                (mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_read),        //                                               .read
		.pll_reconfig_0_mgmt_avalon_slave_readdata            (mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_readdata),    //                                               .readdata
		.pll_reconfig_0_mgmt_avalon_slave_writedata           (mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_writedata),   //                                               .writedata
		.pll_reconfig_0_mgmt_avalon_slave_waitrequest         (mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_waitrequest)  //                                               .waitrequest
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
